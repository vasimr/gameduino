
module RAM_SPRIMG (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [14:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [14:0] addrb
    );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB(dib[0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[0]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB(dib[1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[1]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram2 (
      .DIA(dia[2]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[2]),
      .SSRA(ssra),

      .DIB(dib[2]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[2]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram3 (
      .DIA(dia[3]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[3]),
      .SSRA(ssra),

      .DIB(dib[3]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[3]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram4 (
      .DIA(dia[4]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4]),
      .SSRA(ssra),

      .DIB(dib[4]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram5 (
      .DIA(dia[5]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[5]),
      .SSRA(ssra),

      .DIB(dib[5]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[5]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
         .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram6 (
      .DIA(dia[6]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[6]),
      .SSRA(ssra),

      .DIB(dib[6]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[6]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
            .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram7 (
      .DIA(dia[7]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[7]),
      .SSRA(ssra),

      .DIB(dib[7]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[7]),
      .SSRB(ssrb)
      );

endmodule


module RAM_PICTURE (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [12:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [12:0] addrb
    );

    RAMB16_S4_S4 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram0 (
      .DIA(dia[4*0+3:4*0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*0+3:4*0]),
      .SSRA(ssra),

      .DIB(dib[4*0+3:4*0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*0+3:4*0]),
      .SSRB(ssrb)
      );

    RAMB16_S4_S4 #(
          .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram1 (
      .DIA(dia[4*1+3:4*1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*1+3:4*1]),
      .SSRA(ssra),

      .DIB(dib[4*1+3:4*1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*1+3:4*1]),
      .SSRB(ssrb)
      );

endmodule


module RAM_CHR (
    input [1:0] dia, 	// NC
    output [1:0] doa, 	// CHAROUT
    input wea, 		// 0
    input ena,   	// 1
    input clka,		// vga_clk
    input ssra,		// 0
    input [14:0] addra,	// {glyph, row[2:0], _column[2], ~_column[1:0]}
    input [7:0] dib,	// mem_data_wr
    output [7:0] dob,	// mem_data_rd1
    input web,		// mem_wr
    input enb,		// en_chr
    input clkb,		// mem_clk
    input ssrb,		// 0
    input [12:0] addrb	// mem_addr
    );

// 32 across
// Address mode:  AAAAAA / B BBBB, where A is the INIT_A, and B is the bit across the line
//      Note bit 255 .... bit 0
// Note that ASCII 64, hex 0x40 starts at address 0x0400 
    RAMB16_S1_S4 #(
.INIT_00(256'h00C36606060666C3_00C76666C76666C7_00666666E766C381_00C32606E6E666C3),
.INIT_01(256'h00C36666E60666C3_00060606870606E7_00E70606870606E7_0087C6666666C687),
.INIT_02(256'h0066C6870787C666_0083C6C0C0C0C0E1_00C38181818181C3_00666666E7666666),
.INIT_03(256'h00C36666666666C3_006666E6E7E76766_00363636B6F77736_00E7060606060606),
.INIT_04(256'h00C36660C30666C3_0066C687C76666C7_00E0C366666666C3_00060606C76666C7),
.INIT_05(256'h003677F7B6363636_0081C36666666666_00C3666666666666_00818181818181E7),
.INIT_06(256'h00C30303030303C3_00E7060381C060E7_00818181C3666666_006666C381C36666),
.INIT_07(256'h000103F7F7030100_81818181E7C38100_00C3C0C0C0C0C0C3_00CF2603C70321C0),
// Hex 0x20 below
.INIT_08(256'h006666FF66FF6666_0000000000666666_0081000081818181_0000000000000000),
.INIT_09(256'h000000000081C060_00F3667683C366C3_0064660381C06626_0081C760C306E381),
.INIT_0A(256'h00008181E7818100_000066C3FFC36600_000381C0C0C08103_00C08103030381C0),
.INIT_0B(256'h00060381C0603000_0081810000000000_00000000E7000000_0381810000000000),
.INIT_0C(256'h00C36660C16066C3_00E70603C06066C3_00E7818181838181_00C3666667E666C3),
.INIT_0D(256'h0081818181C066E7_00C36666C70666C3_00C3666060C706E7_006060F766E1E060),
.INIT_0E(256'h0381810000810000_0000810000810000_00C36660E36666C3_00C36666C36666C3),
.INIT_0F(256'h00810081C06066C3_000781C060C08107_000000E700E70000_00E08103060381E0),
//       Character 0x40 starts on the line below
.INIT_10(256'h000000FFFF000000_8181818181818181_00E3C1F7F7E3C180_000000FFFF000000),
.INIT_11(256'h0303030303030303_0000FFFF00000000_0000000000FFFF00_00000000FFFF0000),
.INIT_12(256'h0000000E0F838181_00000070F0C18181_8181830F0E000000_C0C0C0C0C0C0C0C0),
.INIT_13(256'h0C0C0C0C0C0CFFFF_0C0E0783C1E07030_3070E0C183070E0C_FFFF0C0C0C0C0C0C),
.INIT_14(256'h0080C1E3F7F7F763_00FFFF0000000000_00C3E7E7E7E7C300_303030303030FFFF),
.INIT_15(256'h00C3E76666E7C300_3C7EE7C3C3E77E3C_8181C1F070000000_0606060606060606),
.INIT_16(256'h818181FFFF818181_0080C1E3F7E3C180_6060606060606060_00C3818166668181),
.INIT_17(256'h103070F0F1F3F7FF_00636367E3300000_8181818181818181_03030C0C03030C0C),
.INIT_18(256'h00000000000000FF_FFFFFFFF00000000_0F0F0F0F0F0F0F0F_0000000000000000),
.INIT_19(256'h3030303030303030_3333CCCC3333CCCC_0C0C0C0C0C0C0C0C_FF00000000000000),
.INIT_1A(256'h818181F1F1818181_3030303030303030_080C0E0F8FCFEFFF_3333CCCC00000000),
.INIT_1B(256'hFFFF000000000000_8181818F8F000000_000000F1F1818181_F0F0F0F000000000),
.INIT_1C(256'h8181818F8F818181_818181FFFF000000_000000FFFF818181_818181F1F1000000),
.INIT_1D(256'h000000000000FFFF_7070707070707070_0E0E0E0E0E0E0E0E_0C0C0C0C0C0C0C0C),
.INIT_1E(256'h0F0F0F0F00000000_FFFF303030303030_FFFFFF0000000000_0000000000FFFFFF),
.INIT_1F(256'hF0F0F0F00F0F0F0F_000000000F0F0F0F_0000008F8F818181_00000000F0F0F0F0),
.INIT_20(256'hFF3C99F9F9F9993C_FF38999938999938_FF99999918993C7E_FF3C99F91919993C),
.INIT_21(256'hFF3C999919F9993C_FFF9F9F978F9F918_FF18F9F978F9F918_FF78399999993978),
.INIT_22(256'hFF993978F8783999_FF7C393F3F3F3F1E_FF3C7E7E7E7E7E3C_FF99999918999999),
.INIT_23(256'hFF3C99999999993C_FF99991918189899_FFC9C9C9490888C9_FF18F9F9F9F9F9F9),
.INIT_24(256'hFF3C999F3CF9993C_FF99397838999938_FF1F3C999999993C_FFF9F9F938999938),
.INIT_25(256'hFFC9880849C9C9C9_FF7E3C9999999999_FF3C999999999999_FF7E7E7E7E7E7E18),
.INIT_26(256'hFF3CFCFCFCFCFC3C_FF18F9FC7E3F9F18_FF7E7E7E3C999999_FF99993C7E3C9999),
.INIT_27(256'hFFFEFC0808FCFEFF_7E7E7E7E183C7EFF_FF3C3F3F3F3F3F3C_FF30D9FC38FCDE3F),
.INIT_28(256'hFF99990099009999_FFFFFFFFFF999999_FF7EFFFF7E7E7E7E_FFFFFFFFFFFFFFFF),
.INIT_29(256'hFFFFFFFFFF7E3F9F_FF0C99897C3C993C_FF9B99FC7E3F99D9_FF7E389F3CF91C7E),
.INIT_2A(256'hFFFF7E7E187E7EFF_FFFF993C003C99FF_FFFC7E3F3F3F7EFC_FF3F7EFCFCFC7E3F),
.INIT_2B(256'hFFF9FC7E3F9FCFFF_FF7E7EFFFFFFFFFF_FFFFFFFF18FFFFFF_FC7E7EFFFFFFFFFF),
.INIT_2C(256'hFF3C999F3E9F993C_FF18F9FC3F9F993C_FF187E7E7E7C7E7E_FF3C99999819993C),
.INIT_2D(256'hFF7E7E7E7E3F9918_FF3C999938F9993C_FF3C999F9F38F918_FF9F9F08991E1F9F),
.INIT_2E(256'hFC7E7EFFFF7EFFFF_FFFF7EFFFF7EFFFF_FF3C999F1C99993C_FF3C99993C99993C),
.INIT_2F(256'hFF7EFF7E3F9F993C_FFF87E3F9F3F7EF8_FFFFFF18FF18FFFF_FF1F7EFCF9FC7E1F),
.INIT_30(256'hFFFFFF0000FFFFFF_7E7E7E7E7E7E7E7E_FF1C3E08081C3E7F_FFFFFF0000FFFFFF),
.INIT_31(256'hFCFCFCFCFCFCFCFC_FFFF0000FFFFFFFF_FFFFFFFFFF0000FF_FFFFFFFF0000FFFF),
.INIT_32(256'hFFFFFFF1F07C7E7E_FFFFFF8F0F3E7E7E_7E7E7CF0F1FFFFFF_3F3F3F3F3F3F3F3F),
.INIT_33(256'hF3F3F3F3F3F30000_F3F1F87C3E1F8FCF_CF8F1F3E7CF8F1F3_0000F3F3F3F3F3F3),
.INIT_34(256'hFF7F3E1C0808089C_FF0000FFFFFFFFFF_FF3C181818183CFF_CFCFCFCFCFCF0000),
.INIT_35(256'hFF3C189999183CFF_C381183C3C1881C3_7E7E3E0F8FFFFFFF_F9F9F9F9F9F9F9F9),
.INIT_36(256'h7E7E7E00007E7E7E_FF7F3E1C081C3E7F_9F9F9F9F9F9F9F9F_FF3C7E7E99997E7E),
.INIT_37(256'hEFCF8F0F0E0C0800_FF9C9C981CCFFFFF_7E7E7E7E7E7E7E7E_FCFCF3F3FCFCF3F3),
.INIT_38(256'hFFFFFFFFFFFFFF00_00000000FFFFFFFF_F0F0F0F0F0F0F0F0_FFFFFFFFFFFFFFFF),
.INIT_39(256'hCFCFCFCFCFCFCFCF_CCCC3333CCCC3333_F3F3F3F3F3F3F3F3_00FFFFFFFFFFFFFF),
.INIT_3A(256'h7E7E7E0E0E7E7E7E_CFCFCFCFCFCFCFCF_F7F3F1F070301000_CCCC3333FFFFFFFF),
.INIT_3B(256'h0000FFFFFFFFFFFF_7E7E7E7070FFFFFF_FFFFFF0E0E7E7E7E_0F0F0F0FFFFFFFFF),
.INIT_3C(256'h7E7E7E70707E7E7E_7E7E7E0000FFFFFF_FFFFFF00007E7E7E_7E7E7E0E0EFFFFFF),
.INIT_3D(256'hFFFFFFFFFFFF0000_8F8F8F8F8F8F8F8F_F1F1F1F1F1F1F1F1_F3F3F3F3F3F3F3F3),
.INIT_3E(256'hF0F0F0F0FFFFFFFF_0000CFCFCFCFCFCF_000000FFFFFFFFFF_FFFFFFFFFF000000),
.INIT_3F(256'h0F0F0F0FF0F0F0F0_FFFFFFFFF0F0F0F0_FFFFFF70707E7E7E_FFFFFFFF0F0F0F0F)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB({dib[6+0],dib[4+0],dib[2+0],dib[0+0]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+0],dob[4+0],dob[2+0],dob[0+0]}),
      .SSRB(ssrb)
      );

    // note: for [A | B] 6C produces [B | A]

    RAMB16_S1_S4 #(
.INIT_00(256'h00C36606060666C3_00C76666C76666C7_00666666E766C381_00C32606E6E666C3),
.INIT_01(256'h00C36666E60666C3_00060606870606E7_00E70606870606E7_0087C6666666C687),
.INIT_02(256'h0066C6870787C666_0083C6C0C0C0C0E1_00C38181818181C3_00666666E7666666),
.INIT_03(256'h00C36666666666C3_006666E6E7E76766_00363636B6F77736_00E7060606060606),
.INIT_04(256'h00C36660C30666C3_0066C687C76666C7_00E0C366666666C3_00060606C76666C7),
.INIT_05(256'h003677F7B6363636_0081C36666666666_00C3666666666666_00818181818181E7),
.INIT_06(256'h00C30303030303C3_00E7060381C060E7_00818181C3666666_006666C381C36666),
.INIT_07(256'h000103F7F7030100_81818181E7C38100_00C3C0C0C0C0C0C3_00CF2603C70321C0),
// Hex 0x20 below
.INIT_08(256'h006666FF66FF6666_0000000000666666_0081000081818181_0000000000000000),
.INIT_09(256'h000000000081C060_00F3667683C366C3_0064660381C06626_0081C760C306E381),
.INIT_0A(256'h00008181E7818100_000066C3FFC36600_000381C0C0C08103_00C08103030381C0),
.INIT_0B(256'h00060381C0603000_0081810000000000_00000000E7000000_0381810000000000),
.INIT_0C(256'h00C36660C16066C3_00E70603C06066C3_00E7818181838181_00C3666667E666C3),
.INIT_0D(256'h0081818181C066E7_00C36666C70666C3_00C3666060C706E7_006060F766E1E060),
.INIT_0E(256'h0381810000810000_0000810000810000_00C36660E36666C3_00C36666C36666C3),
.INIT_0F(256'h00810081C06066C3_000781C060C08107_000000E700E70000_00E08103060381E0),
//       Character 0x40 starts on the line below
.INIT_10(256'h000000FFFF000000_8181818181818181_00E3C1F7F7E3C180_000000FFFF000000),
.INIT_11(256'h0303030303030303_0000FFFF00000000_0000000000FFFF00_00000000FFFF0000),
.INIT_12(256'h0000000E0F838181_00000070F0C18181_8181830F0E000000_C0C0C0C0C0C0C0C0),
.INIT_13(256'h0C0C0C0C0C0CFFFF_0C0E0783C1E07030_3070E0C183070E0C_FFFF0C0C0C0C0C0C),
.INIT_14(256'h0080C1E3F7F7F763_00FFFF0000000000_00C3E7E7E7E7C300_303030303030FFFF),
.INIT_15(256'h00C3E76666E7C300_3C7EE7C3C3E77E3C_8181C1F070000000_0606060606060606),
.INIT_16(256'h818181FFFF818181_0080C1E3F7E3C180_6060606060606060_00C3818166668181),
.INIT_17(256'h103070F0F1F3F7FF_00636367E3300000_8181818181818181_03030C0C03030C0C),
.INIT_18(256'h00000000000000FF_FFFFFFFF00000000_0F0F0F0F0F0F0F0F_0000000000000000),
.INIT_19(256'h3030303030303030_3333CCCC3333CCCC_0C0C0C0C0C0C0C0C_FF00000000000000),
.INIT_1A(256'h818181F1F1818181_3030303030303030_080C0E0F8FCFEFFF_3333CCCC00000000),
.INIT_1B(256'hFFFF000000000000_8181818F8F000000_000000F1F1818181_F0F0F0F000000000),
.INIT_1C(256'h8181818F8F818181_818181FFFF000000_000000FFFF818181_818181F1F1000000),
.INIT_1D(256'h000000000000FFFF_7070707070707070_0E0E0E0E0E0E0E0E_0C0C0C0C0C0C0C0C),
.INIT_1E(256'h0F0F0F0F00000000_FFFF303030303030_FFFFFF0000000000_0000000000FFFFFF),
.INIT_1F(256'hF0F0F0F00F0F0F0F_000000000F0F0F0F_0000008F8F818181_00000000F0F0F0F0),
.INIT_20(256'hFF3C99F9F9F9993C_FF38999938999938_FF99999918993C7E_FF3C99F91919993C),
.INIT_21(256'hFF3C999919F9993C_FFF9F9F978F9F918_FF18F9F978F9F918_FF78399999993978),
.INIT_22(256'hFF993978F8783999_FF7C393F3F3F3F1E_FF3C7E7E7E7E7E3C_FF99999918999999),
.INIT_23(256'hFF3C99999999993C_FF99991918189899_FFC9C9C9490888C9_FF18F9F9F9F9F9F9),
.INIT_24(256'hFF3C999F3CF9993C_FF99397838999938_FF1F3C999999993C_FFF9F9F938999938),
.INIT_25(256'hFFC9880849C9C9C9_FF7E3C9999999999_FF3C999999999999_FF7E7E7E7E7E7E18),
.INIT_26(256'hFF3CFCFCFCFCFC3C_FF18F9FC7E3F9F18_FF7E7E7E3C999999_FF99993C7E3C9999),
.INIT_27(256'hFFFEFC0808FCFEFF_7E7E7E7E183C7EFF_FF3C3F3F3F3F3F3C_FF30D9FC38FCDE3F),
.INIT_28(256'hFF99990099009999_FFFFFFFFFF999999_FF7EFFFF7E7E7E7E_FFFFFFFFFFFFFFFF),
.INIT_29(256'hFFFFFFFFFF7E3F9F_FF0C99897C3C993C_FF9B99FC7E3F99D9_FF7E389F3CF91C7E),
.INIT_2A(256'hFFFF7E7E187E7EFF_FFFF993C003C99FF_FFFC7E3F3F3F7EFC_FF3F7EFCFCFC7E3F),
.INIT_2B(256'hFFF9FC7E3F9FCFFF_FF7E7EFFFFFFFFFF_FFFFFFFF18FFFFFF_FC7E7EFFFFFFFFFF),
.INIT_2C(256'hFF3C999F3E9F993C_FF18F9FC3F9F993C_FF187E7E7E7C7E7E_FF3C99999819993C),
.INIT_2D(256'hFF7E7E7E7E3F9918_FF3C999938F9993C_FF3C999F9F38F918_FF9F9F08991E1F9F),
.INIT_2E(256'hFC7E7EFFFF7EFFFF_FFFF7EFFFF7EFFFF_FF3C999F1C99993C_FF3C99993C99993C),
.INIT_2F(256'hFF7EFF7E3F9F993C_FFF87E3F9F3F7EF8_FFFFFF18FF18FFFF_FF1F7EFCF9FC7E1F),
.INIT_30(256'hFFFFFF0000FFFFFF_7E7E7E7E7E7E7E7E_FF1C3E08081C3E7F_FFFFFF0000FFFFFF),
.INIT_31(256'hFCFCFCFCFCFCFCFC_FFFF0000FFFFFFFF_FFFFFFFFFF0000FF_FFFFFFFF0000FFFF),
.INIT_32(256'hFFFFFFF1F07C7E7E_FFFFFF8F0F3E7E7E_7E7E7CF0F1FFFFFF_3F3F3F3F3F3F3F3F),
.INIT_33(256'hF3F3F3F3F3F30000_F3F1F87C3E1F8FCF_CF8F1F3E7CF8F1F3_0000F3F3F3F3F3F3),
.INIT_34(256'hFF7F3E1C0808089C_FF0000FFFFFFFFFF_FF3C181818183CFF_CFCFCFCFCFCF0000),
.INIT_35(256'hFF3C189999183CFF_C381183C3C1881C3_7E7E3E0F8FFFFFFF_F9F9F9F9F9F9F9F9),
.INIT_36(256'h7E7E7E00007E7E7E_FF7F3E1C081C3E7F_9F9F9F9F9F9F9F9F_FF3C7E7E99997E7E),
.INIT_37(256'hEFCF8F0F0E0C0800_FF9C9C981CCFFFFF_7E7E7E7E7E7E7E7E_FCFCF3F3FCFCF3F3),
.INIT_38(256'hFFFFFFFFFFFFFF00_00000000FFFFFFFF_F0F0F0F0F0F0F0F0_FFFFFFFFFFFFFFFF),
.INIT_39(256'hCFCFCFCFCFCFCFCF_CCCC3333CCCC3333_F3F3F3F3F3F3F3F3_00FFFFFFFFFFFFFF),
.INIT_3A(256'h7E7E7E0E0E7E7E7E_CFCFCFCFCFCFCFCF_F7F3F1F070301000_CCCC3333FFFFFFFF),
.INIT_3B(256'h0000FFFFFFFFFFFF_7E7E7E7070FFFFFF_FFFFFF0E0E7E7E7E_0F0F0F0FFFFFFFFF),
.INIT_3C(256'h7E7E7E70707E7E7E_7E7E7E0000FFFFFF_FFFFFF00007E7E7E_7E7E7E0E0EFFFFFF),
.INIT_3D(256'hFFFFFFFFFFFF0000_8F8F8F8F8F8F8F8F_F1F1F1F1F1F1F1F1_F3F3F3F3F3F3F3F3),
.INIT_3E(256'hF0F0F0F0FFFFFFFF_0000CFCFCFCFCFCF_000000FFFFFFFFFF_FFFFFFFFFF000000),
.INIT_3F(256'h0F0F0F0FF0F0F0F0_FFFFFFFFF0F0F0F0_FFFFFF70707E7E7E_FFFFFFFF0F0F0F0F)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB({dib[6+1],dib[4+1],dib[2+1],dib[0+1]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+1],dob[4+1],dob[2+1],dob[0+1]}),
      .SSRB(ssrb)
      );

endmodule


module RAM_PAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );

    RAMB16_S9_S18 #(
      	.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_SPRVAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [31:0] DIB,
    output [31:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [8:0] ADDRB
    );

    RAMB16_S9_S36 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_SPRPAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );

    RAMB16_S9_S18 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_CODEL (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
  output reg [7:0] ao,
  output reg [7:0] bo
  );
  wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end

      mRAM128X1D
      #( .INIT(0) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
      #( .INIT(0) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
      #( .INIT(0) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
      #( .INIT(0) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
      #( .INIT(0) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
      #( .INIT(0) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
      #( .INIT(0) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
      #( .INIT(0) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));

endmodule


module RAM_CODEH (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
  output reg [7:0] ao,
  output reg [7:0] bo
  );
  wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end

      mRAM128X1D
           #( .INIT(0) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
           #( .INIT(0) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
           #( .INIT(0) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
           #( .INIT(0) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
           #( .INIT(0) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
            #( .INIT(0) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
          #( .INIT(0) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
            #( .INIT(0) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));

endmodule

