
module RAM_SPRIMG (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [14:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [14:0] addrb
    );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB(dib[0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[0]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB(dib[1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[1]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram2 (
      .DIA(dia[2]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[2]),
      .SSRA(ssra),

      .DIB(dib[2]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[2]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram3 (
      .DIA(dia[3]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[3]),
      .SSRA(ssra),

      .DIB(dib[3]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[3]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram4 (
      .DIA(dia[4]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4]),
      .SSRA(ssra),

      .DIB(dib[4]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram5 (
      .DIA(dia[5]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[5]),
      .SSRA(ssra),

      .DIB(dib[5]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[5]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
         .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram6 (
      .DIA(dia[6]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[6]),
      .SSRA(ssra),

      .DIB(dib[6]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[6]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
            .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram7 (
      .DIA(dia[7]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[7]),
      .SSRA(ssra),

      .DIB(dib[7]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[7]),
      .SSRB(ssrb)
      );

endmodule


module RAM_PICTURE (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [12:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [12:0] addrb
    );

    RAMB16_S4_S4 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram0 (
      .DIA(dia[4*0+3:4*0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*0+3:4*0]),
      .SSRA(ssra),

      .DIB(dib[4*0+3:4*0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*0+3:4*0]),
      .SSRB(ssrb)
      );

    RAMB16_S4_S4 #(
          .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram1 (
      .DIA(dia[4*1+3:4*1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*1+3:4*1]),
      .SSRA(ssra),

      .DIB(dib[4*1+3:4*1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*1+3:4*1]),
      .SSRB(ssrb)
      );

endmodule


module RAM_CHR (
    input [1:0] dia, 	// NC
    output [1:0] doa, 	// CHAROUT
    input wea, 		// 0
    input ena,   	// 1
    input clka,		// vga_clk
    input ssra,		// 0
    input [14:0] addra,	// {glyph, row[2:0], _column[2], ~_column[1:0]}
    input [7:0] dib,	// mem_data_wr
    output [7:0] dob,	// mem_data_rd1
    input web,		// mem_wr
    input enb,		// en_chr
    input clkb,		// mem_clk
    input ssrb,		// 0
    input [12:0] addrb	// mem_addr
    );

// 32 across
// Address mode:  AAAAAA / B BBBB, where A is the INIT_A, and B is the bit across the line
//      Note bit 255 .... bit 0
// Note that ASCII 64, hex 0x40 starts at address 0x0400 
    RAMB16_S1_S4 #(
.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
//       Character 0x40 starts on the line below
.INIT_10(256'h07C06306060666C603C06766C66766C607606666E667C68301C02306E6E666C6),
.INIT_11(256'h7711D37777F71777D311171717971717F711F71717971717F71197D7777777D7),
.INIT_12(256'h7171177D7971797D7771193D7D1D1D1D1F111D39191919191D311777777F7777),
.INIT_13(256'h77D711D37777777777D3117777F7F7F7777711373737B7F7773711F717171717),
.INIT_14(256'h191F711D37771D31777D31177D797D77777D711F1D377777777D311171717D77),
.INIT_15(256'hD37777113777F7B73737371191D3777777777711D37777777777771191919191),
.INIT_16(256'h71331D111D31313131313D311F7171391D171F711919191D3777777117777D39),
.INIT_17(256'h11111111111113F7F713111191919191F7D3911111D3D1D1D1D1D1D311DF3713),
.INIT_18(256'h1D317F391117777FF77FF7777111111111177777711911111919191911111111),
.INIT_19(256'h13131391D1111111111191D17111F3777793D377D31175771391D177371191D7),
.INIT_1A(256'h1111111111111119191F7919111111177D3FFD37711111391D1D1D1911311D19),
.INIT_1B(256'h777777F777D311171391D1713111119191111111111111111111F71111111391),
.INIT_1C(256'h171F777F1F17111D37771D17177D311F71713D17177D311F791919193919111D),
.INIT_1D(256'hD37777D37777D31191919191D177F711D37777D71777D311D3777171D717F711),
.INIT_1E(256'h1F19113171391F11391911111911111111191111191111111D37771F37777D31),
.INIT_1F(256'h111111FFFF11111111911191D17177D3111791D171D19117111111F711F71111),
.INIT_20(256'h111111111FFFF1111111111FFFF111111919191919191919111F3D1F7F7F3D19),
.INIT_21(256'h11D1D1D1D1D1D1D1D113131313131313131111FFFF111111111111111111FFFF),
.INIT_22(256'hF1DFFFF1D1D1D1D1D1D1111111F1F93919111111171F1D191919191931F1F111),
.INIT_23(256'hD311313131313131FFFF1D1D1D1D1D1DFFFF1D1F1793D1F171313171F1D19317),
.INIT_24(256'h1111117171717171717171191D1F3F7F7F77311FFFF111111111111D3F7F7F7F),
.INIT_25(256'h71717111D391917777919111D3F77777F7D3113D7FF7D3D3F77F3D9191D1F171),
.INIT_26(256'h191919113131D1D13131D1D919191FFFF9191911191D1F3F7F3D191717171717),
.INIT_27(256'h1F1F1F1F1111111111111111113171F1F1F3F7FF11737377F331111191919191),
.INIT_28(256'hD1D1D1D1DFF1111111111111111111111111111FFFFFFFFFF111111111F1F1F1),
.INIT_29(256'h1F9FDFFFFF3333DDDD1111111131313131313131313333DDDD3333DDDD1D1D1D),
.INIT_2A(256'h1F1F1919191F1F1F1F111111111919191F1F19191913131313131313131191D1),
.INIT_2B(256'h11FFFF919191919191F1F1111111FFFF1111111111119191919F9F1111111111),
.INIT_2C(256'hF1F1F1F1F1F1F1D1D1D1D1D1D1D1D9191919F9F919191919191FFFF111111111),
.INIT_2D(256'hFFFF11111111111111111111FFFFFF111111111111FFFF71717171717171711F),
.INIT_2E(256'h111119F9F91919111111111F1F1F1F11F1F1F1F11111111FFFF313131313131F),
.INIT_2F(256'hFF99999919993D7FFF3D99F91919993DF1F1F1F11F1F1F1F111111111F1F1F1F),
.INIT_30(256'h9FF19F9F979F9F919FF79399999993979FF3D99F9F9F9993DFF3999993999993),
.INIT_31(256'h1FFF3D7F7F7F7F7F3DFF99999919999999FF3D999919F9993DFFF9F9F979F9F9),
.INIT_32(256'h999FFD9D9D9591999D9FF19F9F9F9F9F9F9FF993979F9793999FF7D393F3F3F3),
.INIT_33(256'h9939FF1F3D999999993DFFF9F9F939999939FF3D99999999993DFF9999191919),
.INIT_34(256'h99999FF3D999999999999FF7F7F7F7F7F7F19FF3D999F3DF9993DFF993979399),
.INIT_35(256'h3F9F19FF7F7F7F3D999999FF99993D7F3D9999FFD9991959D9D9D9FF7F3D9999),
.INIT_36(256'h93D7FFFFF3D3F3F3F3F3F3DFF31D9FD39FDDF3FFF3DFDFDFDFDFD3DFF19F9FD7),
.INIT_37(256'hFF999999FF7FFFFF7F7F7F7FFFFFFFFFFFFFFFFFFFFFFD1919FDFFFF7F7F7F7F),
.INIT_38(256'h97D3D993DFF9B99FD7F3F99D9FF7F399F3DF91D7FFF99991199119999FFFFFFF),
.INIT_39(256'h3D113D99FFFFFD7F3F3F3F7FFDFF3F7FFDFDFD7F3FFFFFFFFFFF7F3F9FFF1D99),
.INIT_3A(256'hFFFFFFFFFFFFFFFFFFF19FFFFFFFD7F7FFFFFFFFFFFFFFF7F7F197F7FFFFFFF9),
.INIT_3B(256'hF9FD3F9F993DFF197F7F7F7D7F7FFF3D99999919993DFFF9FD7F3F9FDFFFFF7F),
.INIT_3C(256'hD999939F9993DFF3D999F9F39F919FF9F9F19991F1F9FFF3D999F3F9F993DFF1),
.INIT_3D(256'hFF7FFFFF7FFFFFFF3D999F1D99993DFF3D99993D99993DFF7F7F7F7F3F9919FF),
.INIT_3E(256'hFF97F3F9F3F7FF9FFFFFF19FF19FFFFFF1F7FFDF9FD7F1FFD7F7FFFFF7FFFFFF),
.INIT_3F(256'h7F7F7F7F7F7F7F7FFF1D3F19191D3F7FFFFFFF1111FFFFFFFF7FFF7F3F9F993D)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB({dib[6+0],dib[4+0],dib[2+0],dib[0+0]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+0],dob[4+0],dob[2+0],dob[0+0]}),
      .SSRB(ssrb)
      );

    RAMB16_S1_S4 #(
.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
//       Character 0x40 starts on the line below
.INIT_10(256'h17D17317171777D713D17777D77777D717717777F777D79311D13317F7F777D7),
.INIT_11(256'h6600C36666E60666C300060606870606E700E70606870606E70087C6666666C6),
.INIT_12(256'h6060066C6870787C6660083C6C0C0C0C0E100C38181818181C300666666E7666),
.INIT_13(256'h66C700C36666666666C3006666E6E7E7676600363636B6F7773600E706060606),
.INIT_14(256'h181E700C36660C30666C30066C687C76666C700E0C366666666C300060606C76),
.INIT_15(256'hC36666003677F7B63636360081C3666666666600C36666666666660081818181),
.INIT_16(256'h70321C000C30303030303C300E7060381C060E700818181C3666666006666C38),
.INIT_17(256'h00000000000103F7F703010081818181E7C3810000C3C0C0C0C0C0C300CF2603),
.INIT_18(256'h0C306E381006666FF66FF6666000000000066666600810000818181810000000),
.INIT_19(256'h03030381C0000000000081C06000F3667683C366C30064660381C066260081C7),
.INIT_1A(256'h1000000000000008181E7818100000066C3FFC36600000381C0C0C0810300C08),
.INIT_1B(256'h666667E666C300060381C0603000008181000000000000000000E70000000381),
.INIT_1C(256'h060F766E1E06000C36660C16066C300E70603C06066C300E781818183818100C),
.INIT_1D(256'hC36666C36666C30081818181C066E700C36666C70666C300C3666060C706E700),
.INIT_1E(256'h0E08103060381E00381810000810000000081000081000000C36660E36666C30),
.INIT_1F(256'h000000FFFF00000000810081C06066C3000781C060C08107000000E700E70000),
.INIT_20(256'h000000000FFFF0000000000FFFF000000818181818181818100E3C1F7F7E3C18),
.INIT_21(256'h00C0C0C0C0C0C0C0C003030303030303030000FFFF000000000000000000FFFF),
.INIT_22(256'hE0CFFFF0C0C0C0C0C0C0000000E0F83818100000070F0C181818181830F0E000),
.INIT_23(256'hC300303030303030FFFF0C0C0C0C0C0CFFFF0C0E0783C1E070303070E0C18307),
.INIT_24(256'h0000006060606060606060080C1E3F7F7F76300FFFF000000000000C3E7E7E7E),
.INIT_25(256'h60606000C381816666818100C3E76666E7C3003C7EE7C3C3E77E3C8181C1F070),
.INIT_26(256'h181818103030C0C03030C0C818181FFFF8181810080C1E3F7E3C180606060606),
.INIT_27(256'h0F0F0F0F0000000000000000103070F0F1F3F7FF00636367E330000081818181),
.INIT_28(256'hC0C0C0C0CFF0000000000000000000000000000FFFFFFFFFF000000000F0F0F0),
.INIT_29(256'h0F8FCFEFFF3333CCCC0000000030303030303030303333CCCC3333CCCC0C0C0C),
.INIT_2A(256'h0F1F1818181F0F0F0F000000000818181F1F18181813030303030303030080C0),
.INIT_2B(256'h00FFFF818181818181F1F1000000FFFF0000000000008181818F8F0000000000),
.INIT_2C(256'hE0E0E0E0E0E0E0C0C0C0C0C0C0C0C8181818F8F818181818181FFFF000000000),
.INIT_2D(256'hFFFF00000000000000000000FFFFFF000000000000FFFF70707070707070700E),
.INIT_2E(256'h000008F8F81818100000000F0F0F0F00F0F0F0F00000000FFFF303030303030F),
.INIT_2F(256'hFF99999918993C7EFF3C99F91919993CF0F0F0F00F0F0F0F000000000F0F0F0F),
.INIT_30(256'h8FF18F9F978F9F918FF78399999993978FF3C99F9F9F9993CFF3899993899993),
.INIT_31(256'h1EFF3C7E7E7E7E7E3CFF99999918999999FF3C999919F9993CFFF9F9F978F9F9),
.INIT_32(256'h899FFC9C9C9490888C9FF18F9F9F9F9F9F9FF993978F8783999FF7C393F3F3F3),
.INIT_33(256'h9938FF1F3C999999993CFFF9F9F938999938FF3C99999999993CFF9999191818),
.INIT_34(256'h99999FF3C999999999999FF7E7E7E7E7E7E18FF3C999F3CF9993CFF993978389),
.INIT_35(256'h3F9F18FF7E7E7E3C999999FF99993C7E3C9999FFC9880849C9C9C9FF7E3C9999),
.INIT_36(256'h83C7EFFFF3C3F3F3F3F3F3CFF30D9FC38FCDE3FFF3CFCFCFCFCFC3CFF18F9FC7),
.INIT_37(256'hFF999999FF7EFFFF7E7E7E7EFFFFFFFFFFFFFFFFFFFEFC0808FCFEFF7E7E7E7E),
.INIT_38(256'h97C3C993CFF9B99FC7E3F99D9FF7E389F3CF91C7EFF99990099009999FFFFFFF),
.INIT_39(256'h3C003C99FFFFFC7E3F3F3F7EFCFF3F7EFCFCFC7E3FFFFFFFFFFF7E3F9FFF0C99),
.INIT_3A(256'hEFFFFFFFFFFFFFFFFFF18FFFFFFFC7E7EFFFFFFFFFFFFFF7E7E187E7EFFFFFF9),
.INIT_3B(256'hF9FC3F9F993CFF187E7E7E7C7E7EFF3C99999819993CFFF9FC7E3F9FCFFFFF7E),
.INIT_3C(256'hC999938F9993CFF3C999F9F38F918FF9F9F08991E1F9FFF3C999F3E9F993CFF1),
.INIT_3D(256'hFF7EFFFF7EFFFFFF3C999F1C99993CFF3C99993C99993CFF7E7E7E7E3F9918FF),
.INIT_3E(256'hFF87E3F9F3F7EF8FFFFFF18FF18FFFFFF1F7EFCF9FC7E1FFC7E7EFFFF7EFFFFF),
.INIT_3F(256'h7E7E7E7E7E7E7E7EFF1C3E08081C3E7FFFFFFF0000FFFFFFFF7EFF7E3F9F993C)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB({dib[6+1],dib[4+1],dib[2+1],dib[0+1]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+1],dob[4+1],dob[2+1],dob[0+1]}),
      .SSRB(ssrb)
      );

endmodule


module RAM_PAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );

    RAMB16_S9_S18 #(
      	.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_SPRVAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [31:0] DIB,
    output [31:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [8:0] ADDRB
    );

    RAMB16_S9_S36 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_SPRPAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );

    RAMB16_S9_S18 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_CODEL (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
  output reg [7:0] ao,
  output reg [7:0] bo
  );
  wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end

      mRAM128X1D
      #( .INIT(0) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
      #( .INIT(0) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
      #( .INIT(0) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
      #( .INIT(0) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
      #( .INIT(0) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
      #( .INIT(0) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
      #( .INIT(0) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
      #( .INIT(0) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));

endmodule


module RAM_CODEH (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
  output reg [7:0] ao,
  output reg [7:0] bo
  );
  wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end

      mRAM128X1D
           #( .INIT(0) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
           #( .INIT(0) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
           #( .INIT(0) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
           #( .INIT(0) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
           #( .INIT(0) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
            #( .INIT(0) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
          #( .INIT(0) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
            #( .INIT(0) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));

endmodule

