`define ALTERA
`define GENERIC_RAM

module RAM_SPRIMG (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [14:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [14:0] addrb
    );
`ifdef GENERIC_RAM
	srambDrsws #(
		.DATA_WIDTH(8),
		.ADDR_WIDTH(15)
	) ram (
		.DIA(dia),
      .WEA(wea),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa),

      .DIB(dib),
      .WEB(web),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob),
	);
	
`elsif ALTERA
	RAMB16_S8_S8 ram (
	    .DIA(dia),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa),
      .SSRA(ssra),

      .DIB(dib),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob),
      .SSRB(ssrb)
	);

`else
    RAMB16_S1_S1 #(
      .INIT_00(256'b0000000000010001000000000000000100000000001000110000000000000011000000000000011100000000110001110000000000001111000000010001111100000000001111110000011000111111000011000111111100011000111111110010000111111111010000111111111110000111111111111000111111111111),
.INIT_01(256'b0000000000000100000000000000010000000000000001000000000000000000000000000000001010000000000000101000000000000000000000000000000110000000000000001100000000000000110000000000000110000000000000011000000000000000100000000000000011000000000000001100000000000000),
.INIT_02(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111100111111111111110001111111111111000011111111111100000111111111110000001111111111000000011111111100000001111111111001000011111111),
.INIT_03(256'b0011101000000001011101010000000000111110100000010111111101010000111111111010101111111111110101101111111010101000111111111101000011111110101000001111111111000000111111111010000011111111000000001111111010000000111111110000000011110110000000001110010000000000),
.INIT_04(256'b1111000010000000111110000100000011111000101000001111110000010000111111000000000011111100000000001111110001000010111111000100000011111100010100111111110001101010111111000101010111111100011111111111110001010101111111000111111111111100011111111111110001111111),
.INIT_05(256'b1111111111111111111111111111111101111111111111110001111111111111000001111111111100000001111111110000000011111111100010000011111111100000000011111111000100000111111100001000000111110000000000001001110000010000110101100000100011110101100001001111100101100000),
.INIT_06(256'b1111111111000001111111111000001111111111000001111111110000101111111110000101111111110000101111111100001011111111000001011111111100000111111111110010111111111111101111111111111111111111111111111111111111111111111111111111111111111111111110001111111111101101),
.INIT_07(256'b0111111111111111001111111111111100011111111111111000111111111111010001111111111100000011111111110000000111111111100000001111111101000000011111111110001000111111111110000011111110101100000111111011100000001111101111011100011100111111110000111011111111110001),
.INIT_08(256'b1111111111111100111111111111111011111111111111111111111111111111111111111111111101011111111111111000000011100111010111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_09(256'b0000000101011111001000000010101000100010000000010011101000000001010111111111111100111111111111110101011111111111001111111111111101010111111111111011111111111111010111111111111110111111111111110111111111111111100101111111111111010111111111110000011011000100),
.INIT_0A(256'b1111101000111110011110000000001100001011111111110101010111111111000010101011111100000101011111110000101010111111000001011111111100000010101111110001010111111111000000101111111101010101111111111001111111000101000000000000000000000000000000011111111111111111),
.INIT_0B(256'b0000101111111111000001011111111100001011110101000001011111110000000001111000000000010000000000000000000000001111000000000111111100000011111111110000111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001),
.INIT_0C(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111110000000011111000000000001000000000000110000000001000111100000100111111110100111111111111),
.INIT_0D(256'b1111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111001111111111111100011111111111110000011111111111010000011111111101000000011111110010100000001111001101100000000001110101100000000110101101010000),
.INIT_0E(256'b1111111111000111111111100000111111111111000111111111110000011111111111100011111111111100001111111111101000111111111111000111111111111000011111111111100000000000111111000000000011111000000000001111100000000000111111011111111111111101111111111111111001111111),
.INIT_0F(256'b1111111111111000111111111110000011111111100000011111111100000101111111000001010011111000010100001110000001000000110000100000101010000010000001010001100000001011000100000001011101000000000011111000000000010110000000000000111100000000000011100101000000111010),
.INIT_10(256'b1100000000000000010000000000100001000000000000001100000000011000000000000000100011000000000100010000000000000001100000000000000110000000000000010000000000010001000000000000001100000000000000110000000001000011000000000100011100000000000001100000000001000100),
.INIT_11(256'b0011000110101101111000010001001010000000010010110000000011100011000000001100001100000000000001110000000000101111000000000001011100000000000011110000000000111111000000000011111100000000000011110000000000001111100000000001111110000000000011110000000000011111),
.INIT_12(256'b1000000000000000111000000100000001000000000000001011000000000000010100000000000000100000000000000011000000000000000000000000000000010000000000001001100000000000110000000000000000010100000000010001001000000010000011010000011000000101101010001000000101100000),
.INIT_13(256'b1101001011100000111110100001100011100100000011101111110000001110111011000000000011110101000001111111011011001101111101100000110011111011110100001111101010000000111110000100000011111100100000001111110100000000111111010000000011111110000000001011111010001110),
.INIT_14(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111000000011111111000000001111111000010110111111000000000011111100000100001111100010111000),
.INIT_15(256'b0000001001011111000000100100111100000001000101110000000101100111000000000010111100000001001011110000000100010011000000010000010000000001000101110000000000001110000000000000001000000010000010100000001100000111000000110010001100000001000001110000000000100001),
.INIT_16(256'b1111111111111111111111111111111111111111111111111111000000011111011000000000011100000000000000110000011111000001100000110001100011000111100011001001111111000010011011111111101101001100011101010011010110111110000110101111111100001111011111110000001011111111),
.INIT_17(256'b1000000000000000000000000001000010000000000000000000000000000000000000000000000000001000000000000001000000000000000010000000000000110100000000000001100000000000000111100000000000100100000000000101011000000000000010100000000001000101000000000100001000000000),
.INIT_18(256'b1111111111111111111111111100001111111111100000001111111100000000111111100000110011111100010111011111100001000001111100010111111000110001100111110000001010001100000000101001100001000000110100010011001011010100111010001110100011111000110110000111110111110000),
.INIT_19(256'b1111111111011110111111111111110111111111111111101111111111111101111111111111111011111111111111001111111111111110011111111111110011111111111111100111111111111100011111111111101010111111111111000111111111111000101111111111110100111111111110100111111111111101),
.INIT_1A(256'b1111111111111111111111111111111111111111111111111111111111111111000011111111100000000111111100000000001111100000110100011100011011100000100011100011000010011001000111000000000001011010000101100010101000110110111110000001011011111101110110001111111010111101),
.INIT_1B(256'b0000001111111110011111111111111111111111111111100101111111111110111111111111111101111111111111111111111111111110111111111111111000000111111111100101111111111111110011111111111100100111111111010001111111111110010011111111111100011111111111011101111111111001),
.INIT_1C(256'b0111111111111111001111111111111100011111111111110000111111111111100000111111100011000001111100001001000011100000110001000000010111110100000011101111110100001100111111111100000011111111110110001111111001001100111111111001100011111111101010011111111111111101),
.INIT_1D(256'b0000000011010001000000011100001000000010100001010001001000000011010111000000010101000010000010110011010000000111001010000000101100110100000101100011000000001001000100000010001000001000010101100001000010100010000100010101101000000010110100100000010101010010),
.INIT_1E(256'b1110000010101010111000001000011100000011101010000000001000101111000000010000000001100111100111111011011110111111010110100111111100111000011111111001110001111111000010001111111100000001001111110000000010011111000000000100111100000000001011110000000000010111),
.INIT_1F(256'b0000000000011001000000000000000110000000000100011000000000010001000001010000100100000000000000011001010101000001100000100000100110010101010110011010101010000001001101010111001100111010101000110001111111010011000010101000001100000111100001110011000000001111),
.INIT_20(256'b0000000000010111000000000011111100000000011111110000000000111111000000000011111000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010000000000000011000000001010101),
.INIT_21(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110000110000011000000010000000000000000000000000010110),
.INIT_22(256'b1110010000000000111011000000000011101000000000001110101000000000111010100000000011000111010100001100001010000000110011010101000011000110101000001100010101010100100001111010100110010101010101011000111111111000100101110101010000011111111110010001111111110101),
.INIT_23(256'b0100000100001111110000011100011100001001110000110100001111000001101000111100100001000001011010001010100000100100010000000110010010101000011100000000000000110000000000000000010100000000000001000000000000001001100000000000001101000000000001100010000000000000),
.INIT_24(256'b1111100000000111111110100100011111111100011000111111110101100011111111110001001011111111101000101111111101100010111111111111000011111111111100001111111111100001111111111101000111111111111000000111111101100000001111110010000110011001000000000010110100001000),
.INIT_25(256'b1111111111100110111111111011011011111111011010101111111100000100111111111100100011111111010100001111111010000000111111001010000011111101000000111111111001000111111110010000011111111010100011111111101010001111111101100000111111110010000111111111101100011111),
.INIT_26(256'b1100010110011111001000011000111100011001000001110000100100011111000011010000001100000001000011110000000100000001000000010000000000000011000000110000000110010001000000111001100000000001000111000000011110011110000000010011111100001000001111110100100001111111),
.INIT_27(256'b0000000000000011000000010011000100000000001100110000000100110111000000001010011100000001001000110000000100101111000000011010011100000000101001110000000100001111000000000101011100000000110011110000000011111111000000001111111100000000111011110000000011111111),
.INIT_28(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111000000000111111000000000001111000101011100011100110110000000110011110101010011000111110011000100011011100000010111111100010001),
.INIT_29(256'b0000000000001000000000000000010000000000000011000000000001000000001001000100000000000100010000001010000001001000010101100100100010100101010010000101001011001000101000010100110011110111110000011010111110000000111101111000000010111111100001111111001110000111),
.INIT_2A(256'b1100010011111011101000100111101111010001111101001010000011100010110000000111010010101000111000001100000000010000101010000010010011000000010001001010100000100000110000000100100010100000010010001101000000001000101000000000100011010000000011001000000001001100),
.INIT_2B(256'b1100111111111110010001111111111111001011111111110100011111111111110000011111111111000001111111111100000111111111110000011111111111000001111111110000000001111111001000001011111111000000011111110100001000010010111000110000100111000111100000000000111111000000),
.INIT_2C(256'b0101110000101011111111010101101101011110001111011111111001011101111111100011111111111111111111111111111110111111111111110011111111111111111111111111111110111110111111111001110011111111111111001111111111111110111111111111111011111111110011001111111111101100),
.INIT_2D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111110000111111111111000001111111111100000011111111111101000111111111000110001111111111110000011111111100101000111110000111100011110000101101000110000001111100010001),
.INIT_2E(256'b0100000000000000010000000000000011000000000000000000000000001000010000000000100001000000000010000000000000000000000000000000000000000000000000000000000000001010010000000000100001000000000010100100000000001101010000000000101001000000000011110100000000001101),
.INIT_2F(256'b0000011000000000100001000000000100000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000100000000000010100000000000000101),
.INIT_30(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111100111111111111110001111111111111000011111111111100000111111111111010001111111111010000011111111100100000111111111011010001111111),
.INIT_31(256'b1111111110101001111111111111000111111111101010100111111111110010111111111110100001111111111110001111111100100000111111001000000011111010000001001111000000011100100100000011110010000000111111000000001111111100000011111111110001111111111111001111111111111100),
.INIT_32(256'b0000010110111101000000100111101000000101011111000000101100101010000001110001110010000111000101100000111100010100000011111000100011011111000010000001111000000100000111110000100001011100000000000001111000000000001110000100010011110100010000000011100010001000),
.INIT_33(256'b0000011111111111000000001111111101000000001111111101000000001111000110100000011100000110100000010000000111000000000000000111000000000000001101000000000000001010000000000000011100000000000000110000000000000001000000000000000010000000000000000110000000000100),
.INIT_34(256'b0000000000000011000000000000010100000000000010110000000000000101100000000010101100000000000001011000000000101011000000000000011100000000000011101010000000010110000111111111000010000000000000001100000000000000010000000000111100100000011111110000100000000111),
.INIT_35(256'b0000000000101100000000000000001000000000010110100000000000001101000000000101011000000000000011100000000001010111000000000000101100011000000101110001000000001011101000000000011110000000000010110000001000000111000000100000101100001110000001110100100000001110),
.INIT_36(256'b1000010101001110000010101000000100000111110000000000111110100000010101111101000000101111011010100001011011010000001011100110100001011110111101000011111001111010011100000011111000011110000010111000000010001000010100000011110010000000000000010101000000000000),
.INIT_37(256'b1111110010100000111111110000000011111111111000001111111111111000111111111111011011111111111110011111111111111100111111111111110111111111111111100111111111110101101111111111111000011111111101010000011111111110000000101111111111000000110111111111000000111101),
.INIT_38(256'b1111110110111100111111110111110011111111101101101111111101101011111111101111000011111110111010101111111101010000111111110010000011111111000100001111111110001000111111101000000011111111110011001111111010100000111111110100000101111110101010000111111111010000),
.INIT_39(256'b1111111111111010111111111111111111111111111110101111111111111111111111111111111111111111111110101111111110110010111110101001000011110111000000011111100000000000000000000000000100000000100010110000011100010111001111100010110011111110000101001111110001101000),
.INIT_3A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111000000000111110000000000011100000000001101000000110000111),
.INIT_3B(256'b1111111111111011111111111111110111111111111111111111111111111100101111111111111000011111111111110000111111111111000001111111111100000011111111110000010111111111000000111111111100000001111111110000000111011111000000101110111100000001111001110000000010110011),
.INIT_3C(256'b0000101111111110000001111111101100001011111011000001010110110000000000111100000000000100100000110000100000001111000001110001111100001101000111110000000000111111000110000011111100000010001111110011001000111110000000100011110001001110001111000000110001111000),
.INIT_3D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100001111111111100000111111111000001011111111000010001111111000010001111111000100101111111000100101011111000100101010),
.INIT_3E(256'b1000000000000001100000000000000100000000000000001000000000000000100000000000000110000000000000001000000000000000000000000000000010000000000000000100000000000001000000000000000101000000000000010000000000000011001000000000001000000000000000110010000000000000),
.INIT_3F(256'b1111111111111111111111111111111111111111111111101111111111111100111111111111110011111111111110001111111111110000111111111110000111111111111000011111111111000010111111111000100011111111000100001111111000000000111111100000000011111100000000001111100010000000)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB(dib[0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[0]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(256'b0000000000001111000000000000111100000000000111110000000000011111000000000111111100000000001111110000000001111111000000011111111100000011111111110000000111111111000000111111111100000111111111110000111111111111000111111111111100111111111111110111111111111111),
.INIT_01(256'b0000000000000011000000000000011100000000000000110000000000000001000000000000001100000000000000010000000000000001100000000000000010000000000000001000000000000001100000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000),
.INIT_02(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111001111111111111100011111111111110000111111111111),
.INIT_03(256'b1101101000000001101101010000000010111110100000010111111101010001111111111010101011111111110101001111111010101100111111111101100011111110101100001111111111100000111111111110000011111111100000001111111110000000111111010000000011111010000000001111010000000000),
.INIT_04(256'b1111111110000000111111110100000011111111001000001111111110010000111111111000100011111111100001001111111110000000111111111000001011111111100100101111111110101011111111111001010111111111101111111111111110010101111111111011111111111111101111111111111110111111),
.INIT_05(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111110001111111111111100001111111111111100011111111111111000011111111111100000111111111110000001111110111110000001111110011100000011111110011100000111111100011100001),
.INIT_06(256'b1111111111111101111111111111101111111111111101111111111111001111111111111001111111111111001111111111110011111111111110011111111111110111111111111100111111111111001111111111111111111111111111111111111111111111111111111111111011111111111111011111111111110111),
.INIT_07(256'b1111111111111111111111111111111111111111111111110111111111111111101111111111111111011111111111111110111111111111011101111111111100111011111111110111110111111111000101111111111101111010111111110111110101111111011111110011111111111111100111111111111111001111),
.INIT_08(256'b1111111111111100111111111111111011111111111111111111111111111111111111111111111111111111111111110000000000011111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_09(256'b0000000101011111111000000010101010011110000000011111100111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100111111111111111100011111100),
.INIT_0A(256'b1111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111000011111111111111111111111111111111111111111111111111),
.INIT_0B(256'b1111111111111111111111111111111111111111111100101111111110101111111111010111111111111011111111111110111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0C(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111110000111111111000111111111000111111111111),
.INIT_0D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111011111111111111110011111111111111111011111111111110011011111111100011011001111),
.INIT_0E(256'b0000000010111111000000010111111100000000111111110000001011111111000000011111111100000001111111110000010111111111000001111111111100000011111111110000001111111111000001111111111100000101111111110000011000000000000000011111111100000010111111110000000111111111),
.INIT_0F(256'b1111111111111111111111111111111111111111111111101111111111111001111111111110011111111111100111111111111101111111111111001111010111111011111110101110111111110100110111111110100011111111111100001111111111101000111111111111001011111111111100101111111111010001),
.INIT_10(256'b0100000000001111010000000000111101000000000001111100000000000111100000000001011101000000000111110000000000001111100000000001111110000000000011110000000000101111000000000001111100000000001111110000000000011111000000000111111100000000011111110000000010111111),
.INIT_11(256'b0011011100101110111000100001010110000001100011100000000011001000000000000000110000000000011100000000000000011000000000000000100000000000001000000000000000010000000000000001000000000000000100000000000000010000000000000000000000000000000100001000000000000000),
.INIT_12(256'b0000000000000000000000000000000010100000000000000111000000000000100100000000000011010000000000001101000000000000111000000000000011100000000000001111100000000000011100000000000011011100000000011110101000000011111100010000000011111011000100111111111001101111),
.INIT_13(256'b1100110011100111111100111111101111100111111111111110111111111111111011111111111111110110111110011111111100101001111100110001110011111010101100001111111001000000111110001100000011111111100000001111110100000000111111010000000011111110000000101011111010001110),
.INIT_14(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110111111111101111111111111101011111111111101000111),
.INIT_15(256'b1111111001101111111111101110111111111111101001111111111110111111111111111111011111111111110100111111111111111011111111111110100011111111111010111111111011111000111111101111010111111110111101001111111011111100111111101111100011111100111110001111111111111110),
.INIT_16(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111011111011101001111011110101000011110110111000000111101001100000000011000010000001000011110100101111110111101010111111111111101111111111111110111111111),
.INIT_17(256'b0111111111101111111111111111111101111111111111111111111111111111111111111111111111100111111111111110111111111111111111111111111111110011111111111100011111111111111111011111111111000011111111111100111111111111101100011111111110111111111111111111101011111111),
.INIT_18(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111001111111111100111001111111101111111111111101000000111111111000000001111110100000000111111010001110000111101000100001110110100000011000101110011011100001111001001110000001100001111),
.INIT_19(256'b0000000000100001000000000000001000000000000000010000000000000010000000000000000100000000000000110000000000000001100000000000001110000000000000010000000000000011000000000000010101000000000000111000000000000111110000000000001001000000000001011100000000000010),
.INIT_1A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100000010111111101010000101111100000000001111111000011111101110001100001111111100110000001101110010100000010001000100000000010000000),
.INIT_1B(256'b0000000000000001000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000001010000000000000010000000000000100010000000000100010000000000011001000000000001101000000000000110000000000000101),
.INIT_1C(256'b1111111111111111111111111111111111111111111111111111111111111111011111111111111100011111111111110011111111111111000110111111100100001001111101000000010111111000000000001010100000000001011100010000000100010011000000001011001000000000000110000000000000001100),
.INIT_1D(256'b0000000000100000000000000000000000000001000000000000101100000000111011100000000000100000000000001101000000000000110111000000000011001000000000001100000000000000110010000000001011000000000001001101000000000100110000000000010011000000000111001100000000011100),
.INIT_1E(256'b1111111100111001111111100000001011111100111011011111111011010001111111111100000011101001100000000000110000000000000001000000000000000110000000000100111100000000000001000000000000000000000000000000000001000000000000000010000000000000000100000000000000001000),
.INIT_1F(256'b1000000000011111100000000001111100000000000011111000000000001111000000000000111110000000000001110000000000000111000000000000011100000000000001110000000000011111100000000001111110000000001011111100000000001111001000000101111110001001101111111110000101111111),
.INIT_20(256'b0000000000000000000000000010000000000000000000000000000000000001000000000100000000000000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001),
.INIT_21(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111),
.INIT_22(256'b1111110000000000111101000000000011110100000000001111010000000000111101000000000011110000000000001111010000000000111110000000000011111000000000001111000000000000111110000000000011100000000000001110100000000001111110000000000011100000000000011110000000000000),
.INIT_23(256'b0110000001111111001100000111111100001000000111110000011000101111000000010011011100000000000111110000000010011011000000000101111100000000000011110000000000011101000000000001001000000000000000100000000000000011000000000000000010000000000000111000000000000000),
.INIT_24(256'b0000000000111111000001100111111100000000000111110000001100111111000000010010111100000000000011110000000011001111000000000001111100000000010111110000000001001110000000000110111100000000001111111000000010011111010000010001111101111010011111101100110011111111),
.INIT_25(256'b0000000000011000000000000110111000000000110110000000000000100011000000001000011100000001010011110000000100011111000000101001111100000000001111110000001100111111000001010111111100000000011111110000010001111111000011001111111100001000111111110000100011111111),
.INIT_26(256'b0001010011100000110010001110000011100100111110001111000011100000111101001111110011111100111100001111110011111110111111001111110111111110111111011111111011111110111111001111111111111110011111111111111001111111111111011111111111110011111111111010001111111111),
.INIT_27(256'b1111111100001010111111100000111011111111000010001111111000000000111111110001110011111110100101001111111010011000111111101001100011111111100100001111111000101000111111110011100011111111001100001111111100100000111111110011000011111111001100001111111100100000),
.INIT_28(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011111111011000010111111110000100101111101000110001111111011011000111111011110100001111),
.INIT_29(256'b1111101111111011111110111111101111111011111101111111101111110111111111111111111111111111111101111111111111111111111110011111111111111010111101111111100101110111111110101111011111111100011110011111110000111111111111000011111111111100001110101111100000110001),
.INIT_2A(256'b1111100100001100111111010000111111111110100010111111111100011011111111110000101111111111100110111111111110101111111111111001101111111111111110111111111111011011111111111011101111111111101110111111111110111111111111111011111111111111101111111111111110111111),
.INIT_2B(256'b0111011111111111111101111111111101110111111111111111101111111111011110011111111101111111111111110111111111111111011111001111111101111110111111111111111011111111111111111011111100111111110111110011111111001001001111111111000001111111111111111111111111111111),
.INIT_2C(256'b0101111111111001111111001111100101011110111111111111111111111111111111101111111111111111011111111111111111111111111111110111111111111111101111111111111111111111111111111011111111111111110111111111111111111101111111111101110111111111110111011111111111101101),
.INIT_2D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111101111111111100001011111111110000010111111111000000111111111100000010111111111000000111111110),
.INIT_2E(256'b0000000000000111100000000000011100000000000001111000000000000111110000000000011111000000000001111100000000001111110000000000111111000000000011111100000000001101100000000000111110000000000011011000000000001010100000000000110110000000000010001000000000001010),
.INIT_2F(256'b0000010000000001000001000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000100000000000010100000000000000101),
.INIT_30(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111001111111111111110111111111111111101111111111111111001111111111),
.INIT_31(256'b0000000000000000000000000000000100000000000000111000000000000111000000000000101110000000000001110000000001111111000000010011111100000100111111110001101111111111110011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_32(256'b1111111100000000111111110000000011111111001000001111111101100000111111110111000001111111011100000111111101101000111111110111000000111111111110000011111011110000001111101111010001111101111111000011110111111100001110111111110000110011111111001111011111110100),
.INIT_33(256'b1111111111111111111111111111111100111111111111111100111111111111111110011111111111111110011111111111111110111111111111111110111111111111111100111111111111111001111111111111111011111111111111111111111111111111111111111111111101111111111111111101111111111111),
.INIT_34(256'b1111111111111100111111111111101011111111111101001111111111111010111111111101010011111111111110101111111111010100111111111111100011111111111100010011111111110010111000000000111101111111111111111011111111111111110111111111111111101111111111111111101111111111),
.INIT_35(256'b1111111111000001111111111111010111111111101000101111111111110000111111111010100011111111111100001111111110101000111111111111010011111111111010000100111111110100100111111111100010111111111101000111110111111000111110111111010011101101111110001011111111110001),
.INIT_36(256'b1111101010111110111101010111111111111000001111111111000001011111101010000010111111010000000101011110100000101111110100000001011110100000000010111100000000000101100000011000000100011100010110001111111100001010111111111100000011111111111111101111111111111111),
.INIT_37(256'b1111110111111111111111110111111111111111110111111111111111110111111111111111110111111111111111111111111111111111111111111111111111111111111111110111111111111111011111111111111111001111111111111111001111111111111111101111111111111111100111111111111111010001),
.INIT_38(256'b1111111110111100111111111011110111111111111111111111111101111111111111110111111111111111011111111111111101111111111111111111111111111111101111111111111111011111111111111110111111111111111110111111111111111101111111111111111101111111111111111111111111111111),
.INIT_39(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111100100111111110010111111101101011111111100101111111111100111111111111100111111111111100111111111111100111111111111110110011111111110101111),
.INIT_3A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111000000111),
.INIT_3B(256'b1111111111111111111111111111110111111111111111010111111111111110111111111111111100111111111111110001111111111111000011111111111100000111111111110000011111111111000000101111111100000001011111110000000110111111000000101101111100000001111011110000000010110111),
.INIT_3C(256'b0000101111111110000001111111101000001011111010110001010110101111000000110011111100000101011111110000101011111111000000101111111100000100111111110000100111111111000010011111111100010001111111110001000111111111001000011111111100001101111111110100111111111111),
.INIT_3D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100001111111111100001111111111000101111111111000101011111111000101010),
.INIT_3E(256'b0000000000000000000000000000000000000000000000011000000000000001100000000000000110000000000000001000000000000000000000000000000000000000000000001000000000000001110000000000000111000000000000011000000000000011110000000000001111100000000000001100000000000001),
.INIT_3F(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111110111111111111010011111111111010001111111111110000111111111110000011111111110000001111111110000000)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB(dib[1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[1]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(256'b0000000000001111000000000001111100000000000111110000000000111111000000000011111100000000011111110000000011111111000000001111111100000001111111110000001111111111000001111111111100001111111111110001111111111111001111111111111101111111111111111111111111111111),
.INIT_01(256'b0000000000000111000000000000001100000000000000110000000000000011000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111),
.INIT_03(256'b1110010111111110110010101111111111000001011111101000000010101110000000000101010000000000001010000000000101010000000000000010000000000001010000000000000000000000000000000010000000000000000000000000000010000000000000010000000000000010000000000000010000000000),
.INIT_04(256'b1111111100000000111111111000000011111111110000001111111111100000111111111111000011111111111110001111111111111100111111111111110011111111111011001111111111010100111111111110101011111111110000001111111111101010111111111100000011111111110000001111111111000000),
.INIT_05(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111100011111111111110000111111111111000011111111111100001111111111110000001111111111110000011111111111110000011111111111100000011111),
.INIT_06(256'b1111111111111110111111111111110011111111111110001111111111110000111111111110000011111111110000001111111100000000111111100000000011111000000000001111000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000111),
.INIT_07(256'b1111111111111111111111111111111111111111111111111111111111111111011111111111111100111111111111110001111111111111000011111111111100000111111111110010001111111111011100011111111101111001111111110111110011111111011111110111111101111111101111110111111111011111),
.INIT_08(256'b0000000000000011000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_09(256'b1111111010100000000111111101010110000001111111101111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111100000011),
.INIT_0A(256'b0000000000000000111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111000000111111111111111111111111111111111111111111111111),
.INIT_0B(256'b1111111111111111111111111111111111111111111100011111111110011111111111001111111111110111111111111101111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0C(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111000000001111000000000000),
.INIT_0D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111110001111111111111000000111111111100010000111111110000111000111111),
.INIT_0E(256'b1111111111111111111111111111111111111110111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111011111111111111101111111111111111111111111111111111111111111111110111111111111111000000000011111110000000001111111100000000),
.INIT_0F(256'b1111111111111111111111111111111111111111111111111111111111111110111111111111100011111111111000001111111110000000111111110000000011111100000000001111000000000000111000000000000010000000000000000000000000000000000000000000001000000000000001010000000000011111),
.INIT_10(256'b0011111111110111001111111111011100111111111111111011111111111111111111111111111110111111111111111111111111101111011111111110111101111111111111111111111111111111111111111101111111111111110111111111111111111111111111111111111111111111101111111111111111111111),
.INIT_11(256'b0011000011010000000111101110100101111111011100111111111110110011111111111011011111111111110001111111111111001111111111111100111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_12(256'b0011111111111111001111111111111100111111111111110010111111111111000011111111111100001111111111110000111111111111000111111111111100011111111111110001011111111111100011111111111111101011111111101111010111111101111110101111110111111101111101111111111110011111),
.INIT_13(256'b0011111100011000000011000000010000001000000000000001000000000000000100000000000000000000000000010000100000001110000010000010001100000000100011110000010000111111000001010011111100000010011111110000001011111111000000101111111100000001111111100100000101110101),
.INIT_14(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110000011111111110000001111111110000000),
.INIT_15(256'b0000000110010000000000011000000000000000110010000000000011001000000000001100000000000000111001000000000011100000000000001111001100000000111100100000000111110001000000011111100100000001111110000000000111111000000000011111110000000011111111000000001111111100),
.INIT_16(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110000000111101110000000001110010000000000011000000000000000111000000001111000001000110000001000010010000000000000100000000000000010000000000),
.INIT_17(256'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000011000000000000010100000000000001010000000000000010100000000000011010000000000011110100000000001111010000000000111111100000000),
.INIT_18(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111110000000111111110000000011111110000000001111111000000000111111100001111111111110000110000001111000010000000011100010000000000110001000000000011000100000),
.INIT_19(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000),
.INIT_1A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111100001111111110000000011111110000000000111110000011111011111001100000010111000110000000111100011000000000110000000000000101000100),
.INIT_1B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000010111000000000001010100000000000100000000000000000010000000000000000000000000001001000000000000000000000000000010),
.INIT_1C(256'b1111111111111111111111111111111111111111111111111111111111111111011111111111111101111111111111110000111111111111000001111111111000000011111110000000000011110000000000100111000000000001001000010000000000100010000000000000000000000000010001000000000000100000),
.INIT_1D(256'b0000000001000000000000001000000000000001000000000000011000000000001001100000000011110000000000001110010000000000111010000000000011101000000000001110100000000001111000000000001011100000000001001111000000001000111100000000000011110000000000001111000000010000),
.INIT_1E(256'b1111111111000111111111110000000111111110111011001111110011100000111111011000000000011101000000000000000100000000000000010000000000000001000000000011110100000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F(256'b0000000000000111000000000000011100000000000001111000000000000111100000000000011100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000001111110000000000111110000000000011111100000000111111111010000111111111100000011111111),
.INIT_20(256'b0000000000000000000000000000000000000000000000000000000001000001000000000000001000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100),
.INIT_21(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000),
.INIT_22(256'b1111100000000000111110000000000011111000000000001111100000000000111110000000000011111000000000001111100000000000111100000000000011110000000000001111000000000000111110000000000011111000000000001111000000000000111000000000000111100000000000011111000000000000),
.INIT_23(256'b0110000011111111000100000011111100000000001111110000001000011111000000010000111100000000000001110000000000000111000000000000001100000000001000110000000000010011000000000000000100000000000010010000000000000000000000000000010000000000000000111000000000000011),
.INIT_24(256'b0000010001111111000000100011111100000010001111110000000100011111000000000001111100000000100111110000000001011111000000000100111100000000000011110000000000011111000000000001111000000000010111100000000000111110000000000111111010100110111111111111001111111111),
.INIT_25(256'b0000000000000000000000000010000100000000010001110000000010011111000000001011111100000000001111110000000101111111000000000111111100000010111111110000001011111111000000001111111100000101111111110000010111111111000001011111111100000001111111110000000111111111),
.INIT_26(256'b0000110001110000000000000110000000000100011000000000010001111000000000000111000000000000011111000000000001111000000000000111110000000010011111110000001001111111000000100111111100000010111111110000001011111111000001001111111100001001111111111110011111111111),
.INIT_27(256'b0000000010011100000000001001100000000000100110000000000010011100000000001001000000000000100100000000000010011000000000001001100000000000100110000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000010000),
.INIT_28(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111100000001111111100000100011111110000110000111110011011000011110100001100001111),
.INIT_29(256'b0000000000110000000000000011010000000000001100000000000000110000000001000011100000000100001110000000010000110000000001000011000000000100001110000000010000110000000001000011110000000000001111000000000001111111000000000111111100000000011111000000010001111010),
.INIT_2A(256'b0000000100000110000000000000010000000000100001100000000010000100000000001000000000000000000000000000000000000100000000000000010000000000010001000000000001000100000000000100010000000000010001000000000001000100000000000100010000000000010001000000000001000100),
.INIT_2B(256'b0011000000000000001110000000000000111100000000000011100000000000001111100000000000111110000000000011110000000000001111110000000000111110000000000011111110000000000111110100000000011111101000000001111111101111000111111111111100111111111111110111111111111111),
.INIT_2C(256'b1010001000000110000000100000011010100000000000100000000100000010000000010000001000000000000000100000000010000010000000001000001000000000000000100000000001000010000000000100001000000000000000100000000000100010000000000010001000000000001000100000000000000010),
.INIT_2D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111000011111111111100000111111111110000001111111111000000011111111100000001111111111000000011111111),
.INIT_2E(256'b0011111111111000001111111111100010111111111110001011111111111000111111111111100011111111111110001111111111111000111111111111100011111111111110001111111111111000111111111111100011111111111110001111111111111000111111111111100011111111111110001111111111111000),
.INIT_2F(256'b1111111111111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111101111111111111111011111111111101011111111111111010),
.INIT_30(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111001111111111111100011111111111110000111111111111),
.INIT_31(256'b1111111111111111111111111111111111111111111111101111111111111101111111111111111111111111111011111111111111011111111111110111111111111101111111111111011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_32(256'b0000000001111111000000001011111100000000111111110000000011011111000000001111111100000000111011110000000011111111100000001111011110000000111101111000000111111111100000011111111111000011111111111000001111111111100001111111111110001111111111111000111111111111),
.INIT_33(256'b1111111111111111111111111111111111111111111111110011111111111111000001111111111100000001111111110000000001111111000000000001111100000000000011110000000000000111000000000000000100000000000000000000000000000000000000000000000000000000000000001100000000000000),
.INIT_34(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111110001111111111111111111111111111111110111111111111111001111111111111100011111111111110000011111111111),
.INIT_35(256'b1111111111110100111111111111101011111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111111111011111011111111101111111111111111111111111111111111111011111111111110001111111111100001111111111),
.INIT_36(256'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000011100000001110001111111111110110111111111111111111111111111111111111111111111111),
.INIT_37(256'b1111110000000000111111110000000011111111110000001111111111110000111111111111110011111111111111111111111111111111111111111111111111111111111111110111111111111111101111111111111111101111111111111111101111111111111111001111111111111111000111111111111111100001),
.INIT_38(256'b1111111110000010111111111000001111111111100000011111111100000001111111110000000011111111000000001111111100000000111111111000000011111111100000001111111111000000111111111110000011111111111110001111111111111100111111111111111101111111111111110111111111111111),
.INIT_39(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111100011111111110001111111111100111111111111011111111111111011111111111111001111111111111000111111111111000011111111111000011111111111001111),
.INIT_3A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000),
.INIT_3B(256'b0000000000000011000000000000000100000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000001000000000000000110000000000000101100000000000001111000000000000010110000),
.INIT_3C(256'b0000101111111110000001111111100100001011111001110001010110011111000000110111111100000100111111110000100111111111000000011111111100000011111111110000011111111111000001111111111100001111111111110000111111111111000111111111111100110011111111110011001111111111),
.INIT_3D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111010011111111111010101111111111010101),
.INIT_3E(256'b1000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000001100000000000000110000000000000011000000000000000100000000000000010000000000000001100000000000010110000000000001011000000000000101110000000000001),
.INIT_3F(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111100111111111111100011111111111100001111111111100000111111111100000011111111100000001111111100000000)
    ) ram2 (
      .DIA(dia[2]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[2]),
      .SSRA(ssra),

      .DIB(dib[2]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[2]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_01(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_02(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_03(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111101111111111111101111111111111101111111111111101111111111),
.INIT_04(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_05(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111100001111111111110000011111111111),
.INIT_06(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111000),
.INIT_07(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111100011111111111110000111111111111000001111111111100000001111111110000000011111111000000000111111),
.INIT_08(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_09(256'b1111111111111111111111111111111101111111111111110000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000001111111111111111),
.INIT_0A(256'b1111111111111111000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111111111111111111111111111111111111111111111111),
.INIT_0B(256'b0000000000000000000000000000000000000000000011110000000001111111000000111111111100001111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0C(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111110000111111111),
.INIT_0E(256'b0000000001111111000000001111111100000001111111110000000111111111000000111111111100000011111111110000001111111111000000111111111100000111111111110000011111111111000000111111111100000011111111110000001111111111000000111111111100000001111111110000000011111111),
.INIT_0F(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110001111111111100000),
.INIT_10(256'b1000000000001111100000000000111110000000000011110000000000001111000000000000111100000000000011110000000000011111000000000001111100000000000111110000000000011111000000000011111100000000001111110000000000111111000000000011111100000000011111110000000001111111),
.INIT_11(256'b1100111111111111000000011111111000000000111111000000000001111100000000000111100000000000001110000000000000110000000000000011000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_12(256'b1100000000000000110000000000000011000000000000001100000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111100000000000011110000000000001111100000000000111111000000001111111110000011111111111111111111),
.INIT_13(256'b0001111111111111000111111111111100011111111111110000111111111111000011111111111100001111111111100000011111110000000001111100000000000111000000000000001100000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000011),
.INIT_14(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_15(256'b0000000111100000000000011111000000000001111100000000000111110000000000011111100000000001111110000000000111111100000000011111110000000001111111000000000111111110000000011111111000000001111111110000000111111111000000011111111100000001111111110000000111111111),
.INIT_16(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110000110000111000000000000001100000000000000010000000000000001000000000),
.INIT_17(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000111000000000000011100000000000001111000000000000111100000000000011110000000000),
.INIT_18(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111000001111111111100000111111111100000011111111110000001111111111000000),
.INIT_19(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000),
.INIT_1A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111110010000001111111001000000011111100000000001111111000000000011111000),
.INIT_1B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000011100000000000011100000000000001110000000000000110000000000000111000000000000011),
.INIT_1C(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111110001111111111111000011111111111100000111111111110000001111111111000000011111111100000000111111100000000011111100000000000111110000000000001110000000000000011000),
.INIT_1D(256'b0000000000000000000000000000000000000000000000000000000000000000000110000000000011111100000000001111100000000000111100000000000011110000000000001111000000000000111100000000000111110000000000111110000000000111111000000000111111100000000011111110000000001111),
.INIT_1E(256'b1111111111111111111111111111111111111111000100111111111100000000111111100000000011111110000000001111111000000000111111100000000011111110000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F(256'b1000000000001111100000000000111110000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000111111000000000111111110000000011111111100000011111111111111111111111),
.INIT_20(256'b0000000000001111000000000001111100000000001111110000000000111110000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011),
.INIT_21(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_22(256'b1111100000000000111110000000000011111000000000001111100000000000111110000000000011111000000000001111100000000000111110000000000011111000000000001111100000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001110000000000001),
.INIT_23(256'b1001111111111111000011111111111100000111111111110000000111111111000000001111111100000000111111110000000001111111000000000011111100000000000111110000000000001111000000000000111100000000000001110000000000000111000000000000001110000000000000001100000000000000),
.INIT_24(256'b0000001111111111000000011111111100000001111111110000000011111111000000001111111100000000011111110000000000111111000000000011111100000000001111110000000000111111000000000011111100000000001111110000000001111111100000001111111111000001111111111111111111111111),
.INIT_25(256'b0000000000000000000000000001111000000000001111110000000001111111000000000111111100000000111111110000000011111111000000011111111100000001111111110000000111111111000000111111111100000011111111110000001111111111000000111111111100000111111111110000011111111111),
.INIT_26(256'b0000001111100000000001111111000000000011111100000000001111110000000000111111100000000011111110000000001111111100000000111111111000000001111111100000000111111111000000011111111100000001111111110000000111111111000000111111111100000111111111110001111111111111),
.INIT_27(256'b0000000001111100000000000111110000000000011111000000000001111000000000000111100000000000011110000000000001110000000000000111000000000000011100000000000011110000000000001111000000000000111100000000000011110000000000001110000000000000111000000000000011100000),
.INIT_28(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111001111111111100100111111111000000011111111),
.INIT_29(256'b0000011111111100000001111111100000000111111110000000011111111000000000111111000000000011111100000000001111110000000000111111000000000011111100000000001111111000000000111111100000000011111111100000001111111111000000111111111100000011111111110000001111111100),
.INIT_2A(256'b0000000011111111000000001111111000000000011111000000000001111100000000000111110000000000011111000000000001111000000000000111100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000),
.INIT_2B(256'b1111100000000000111110000000000011111000000000001111110000000000111111000000000011111100000000001111111000000000111111100000000011111111000000001111111100000000111111111000000011111111110000001111111111110000111111111111111111111111111111111111111111111111),
.INIT_2C(256'b0000000111111100000000011111110000000001111111000000000011111100000000001111110000000000111111000000000001111100000000000111110000000000011111000000000000111100000000000011110000000000001111000000000000011100000000000001110000000000000111000000000000011100),
.INIT_2D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111),
.INIT_2E(256'b1100000000000111110000000000011111000000000001111100000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111),
.INIT_2F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_30(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_31(256'b0000000000000000000000000000000000000000000000010000000000000011000000000000011100000000000111110000000000111111000000001111111100000011111111110000111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_32(256'b1111111110000000111111111100000011111111110000001111111111100000111111111110000011111111111100001111111111110000011111111111100001111111111110000111111111111000011111111111100000111111111110000111111111111000011111111111100001111111111110000111111111111000),
.INIT_33(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111),
.INIT_34(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_35(256'b0000000000000011000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111100000000011111110000000001111111000000000111111100000000011111110000000001111110000000000),
.INIT_36(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100000000000001110000000000000001000000000000000000000000000000000000000000000000),
.INIT_37(256'b0000001111111111000000001111111100000000001111110000000000001111000000000000001100000000000000000000000000000000000000000000000000000000000000001000000000000000110000000000000011110000000000001111110000000000111111110000000011111111111000001111111111111110),
.INIT_38(256'b0000000001111111000000000111111000000000011111100000000011111110000000001111111100000000111111110000000011111111000000000111111100000000011111110000000000111111000000000001111100000000000001110000000000000011000000000000000010000000000000001000000000000000),
.INIT_39(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000011111111100001111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110000),
.INIT_3A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_3B(256'b1111111111111100111111111111111011111111111111101111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111011111111111111110111111111111111001111111111111010011111111111110000111111111111101001111),
.INIT_3C(256'b1111010000000001111110000000011111110100000111111110101001111111111111001111111111111011111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_3D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_3E(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111110111111111111111011111111111111110),
.INIT_3F(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111)
    ) ram3 (
      .DIA(dia[3]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[3]),
      .SSRA(ssra),

      .DIB(dib[3]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[3]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(256'b1100000000000000110000000000000011000000000000011100000000000001110000000000000011000000000000011100000000000000100000000000000110000000000000101100000000000000110000000000000010000000000001100000000000000000100000000000000000000000000010000000000000000000),
.INIT_01(256'b0000100001111111000001000111111100100110001111110000001000011111000000010000111100000011100011110000000010000111000000001000001100000000010000110000000000000011000000000000000100000000011000000000000000000000000000000001000000000000000000000000000000010000),
.INIT_02(256'b1100100000000000011101000000000000101000000000000101000000000000111010100000000101010000000000111110101000000010010100000000100010101000001000000100000001100001101010001000011101000011000011111000110000011111010010000111111110000000111111110000001111111111),
.INIT_03(256'b1111110001111111111111000011111111111100001111111111110000111111111111001111111111111000111111111111100001111111111110001111111111110000111111111111000111111111111000110111111111100010001111101100000000010101100011000000101010000000000000010000100000000010),
.INIT_04(256'b1111110000110000111110101000110011111111010000101111101010000010111111110100000111111110100000001111111101000000111111101010000011111101000000001110101010100000110101010000000011110000101000000001000000000000000011000000000000000010000000001100000000000000),
.INIT_05(256'b1111111110011111101111010111111101101011111111111011111111111111111111111111110111111111111111111111111111111101111111111111111111111111111111011111111111111111111111111111110011111111111100101111111110111000111111011100000010011010000000011000000000000111),
.INIT_06(256'b1111111111100001111111111110100111111111111110011111111111110001111111111111100111111111111110011111111111111001111111111110000111111111101000111111111111000111111101110001111110111000011111100000001111111100000111111111110011111111111110001111111111110000),
.INIT_07(256'b1111111111111111111111111111111111010101111111110000000100111111000000000100011100000000000001101111111000000000111111111000000011111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_08(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111000000000001111100000000000000110011111100000000111111000010000011111111100001001111111111110001),
.INIT_09(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111100000111111110000000011110000000000100000000000011011000000001100011100001110000111110000101010111111),
.INIT_0A(256'b1111111111100000111111111100000011111111100000001111111110001001111111111000110011111111100011111111110000000110000000000001011100000000010010110000001011110011000111110011111111110100010110011110100000111111111101000101110011101010001011111111000001010110),
.INIT_0B(256'b0111010111111111000000001011111100000000010111110000001010111111000000000101110110000010100000000100000000000011101000001101000111111111110001111111000100111111010110101111111100010101111111110000101111111111000101010111111100000011111111110001010101111111),
.INIT_0C(256'b1101111111101001001111111111000001111111111011000111111010000011111111110100000011111010100000001111111101010001111110100000000011111111010100010101111010000000000101110101000000000101000000000000000101000000110000000010000011110000001100001111110000000100),
.INIT_0D(256'b1111111101111111111111111111111111111111111010101111111101010000111111111010000011111101010000001111111110101000011111110100000001011111101010000111111111000000000111111110000000001011111100001000001100111010111000000011100011110000000010101111111000000000),
.INIT_0E(256'b1000000000011000010100011000000010000010000000000100000000000000100001000000000000011100000000001011101000000000011101001000000001111010000000001111110101000000111010100000001111111101000010001110101000011100111111010010000011111110110000011111110111000011),
.INIT_0F(256'b0000000010001000000000010100000100000001100000000000000000000100000000000000100000000010000100000000000001000000000100001000000001110000000000011100000110000010100000000000010000001100010010010001111000010011001111110000111101111111100000011111111111000001),
.INIT_10(256'b1000000000011111000000000000111110000000000111110000000000001111000000000001111100000000000011110000000000001111000000000000011100000000000011110000000000001011000000000000001100000000000010010000000000001110010000000000100001000000000010001100000000000000),
.INIT_11(256'b1111111111111110111111111111110011111111111110001111111111110001111111111110000111111111110000101111111110001101111111110001101001111110001101010001111000011110000011000011111100000000111101110110000011111111001100000101011000010000001011110001110100010110),
.INIT_12(256'b1111111100010111101011110000100111111111100110001010111110011100010101111010101010101111111011000001010101001011001010111100110010000101010001111010101011000100000000010100111111000010100011100000000001000111110000001000000011000000010000001010000000000000),
.INIT_13(256'b1111100000111110111110001111000111111000001100111111100000111000111110001101100111111100000001100111110001001110001111000010011000111110001001001001111000000100110111100000001101001110001000011100111000100000100010000001000111000000000100011100000001000001),
.INIT_14(256'b0000000000100011000000100010001100000010001000010000010001100000000000100110000100000000011000000000000001100001000010001110001000001100111000100000000111100001000100011110000000000011111100000011001111110000011001111111000011101111111110000000111111111100),
.INIT_15(256'b0000000011111111000001011111111100000101111111110000000011111111000000001111111100000010011111110000000011111111000000100111111100000001101111110000000101111111000000011011111100000000001111110000000110111111000000100101111100000010101111110000001010111111),
.INIT_16(256'b0100001110000000100000001000000000000000100000000001000011000000000100010000000000010000100000000001000101000000000110001010000000011000000000000011100011100000001110000000000000111100101000000111110001110000011111000000000011111110000000011111111000000100),
.INIT_17(256'b0111000111010000111011011111000000010000010000000000001001110000000001010100000000000000010100000000001100100000000000010010000000000000101100000000000001100000000000001111000001000000010100000000000001100000010000000011000000000000001100000100000000000000),
.INIT_18(256'b0011111111111010011111111111110100111111111110101111111111111110001111111111101110111111111111000111111111111111001111111111110000111111111110000011111111111000001111111111010000011111111110000001111111101001000011111100001100010111111000110001100101000111),
.INIT_19(256'b1111111111011000111111111111111011111111101110001111111100111100111111111010010011111111011011011111111100110010111111111110010111111111101011101111111111111101111111111111111011111111100011011111111111101110111111111101110111111111110111101111111111111101),
.INIT_1A(256'b0011111111111000011111111111000111111111111100011111111111101000111111111111000011111111111000001111111111000000111111111000000011111111010011001111111110011100111111101011110011111111011111101111111011111110111001011111111010010011111111111010011111111111),
.INIT_1B(256'b1111111111101011111111111110010111111111111101111111111111111101101111111111100110111111111111110100111111111101101000111111110101001011111111111000100111111111101001011111111101010000111111110010001011111111000110001111111100001010111111110000011011111111),
.INIT_1C(256'b0000001111010100000001010100000000100011111000010010011101111111000011111111111100000111111111110001101111111111100001111111111110000001111111111100001111111111110001111111111111100000111111111111000101111111111110001001111111111100000110011111111000001011),
.INIT_1D(256'b0000000000001011000000000000000000000000000001110000000000000000000000000000000001000000000000100010000000000001010000000000001110000000000000000000000000000111000000000000000000000000000011100000000000001010000000000000111000000000001001100000000001010010),
.INIT_1E(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000111111000000000001111000000111000),
.INIT_1F(256'b0000000011010000000000000101000010000000000100000000000000010000100000000101000010000000000100000000000001010000100000000001000010000000000100001000000000000000100000000010000010000000000000001000000000100000100000000010100010000000000010001000000000000001),
.INIT_20(256'b0000110010010000001110111010000001000100011000000010011011001111011001101100100011001010111100000100001011000000100000101100000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101),
.INIT_21(256'b0000111111111101001111111111111000111111111110101101111111111100101111111111100011111111111110001111111111111000111111111111010011111111111100010111111111101000111111111111100011111111110100010111111110000001000101100010000100111000010000000000111100000001),
.INIT_22(256'b0110000000000001000100000000001000000000000000010000000000000001100010000000000110000000000000001100000000000001110010000000000011000000000000001100010000000000111001000000000011101100000000001110100000000000111010000000000011101100000000001110110000000000),
.INIT_23(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111100000001111111110000000011111111111000000111111100010000001111110110000000011111),
.INIT_24(256'b1111101100011111111100000001111111110000000111111111000000011111111100100001111111110000000111111111000100011111111100010001111111111001000111111111100000011111111110001000111111110001000011111111100000001111111101000000111111111000010001111111110010000111),
.INIT_25(256'b1111111110000000111111110000000011111110000000011111110000011100111110000011100011110000011001001110000101010000110000110111110110000101111111100000011111110101000011111111111101011111111101010111111111111110101111111111010111111111111110100111111111010000),
.INIT_26(256'b0000000111101111000000011111111100000001111011110000000111101111000000011010111100000001110011110000000000001111000000000000111100000001000011110000011000001111000011100000111110000010000011110000000000001111000001100000111100001100000011111101011010011111),
.INIT_27(256'b1111100100010001100001001001000100000011000100010000000110000001000000010000000100000001000000010000000100000000000000010000000000000001000100000000000101010000000000011001000000000001100100010000000110010001000000010001001100000001000100100000000100000011),
.INIT_28(256'b1111101111001000111111110001000011110011000000001111011000000000111001000000000011111000000000001101101001100000111110000100000010000000001000000000000000100000000001100000000000111110000000001111111100010000111111110001000011111111100010101111111111000000),
.INIT_29(256'b1101000000001000000000000000110001000000110110100000000000011100010000000001111000000000001110000000000111010110000000000011111000000000010111000000001011110110000000111100011000000001111101000000011111100000000001001100001000000001011000100000010010100110),
.INIT_2A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000111111000000000001111100101111100011110110011101000111110011001100001110001000010100000011100010110000100010100110000010011110111100001000100001100001),
.INIT_2B(256'b1111111111000110011111111110111011111111111100000111111111100100101111111111010001111111111111000111111111110000011111111111110000111111111110000101111111111100010111111111100001001111111111010101111111111010011011111111111111000111111110100100011111111111),
.INIT_2C(256'b1011111010000011000111110000001000111111100000111011111101001011000111010000001110111110010101111110110100111111010011101001011001101101001101110011011000011111011001010000101100110110000100100101100000001011101010000000001101011010001010011011110000011001),
.INIT_2D(256'b0100000000001111010000000000111101000000000011110100000000001111010000000000111101000000000011110100000000001110010000000000011000000000000011010100000000001011000000000000000100000000000000110010000000000001001100000000000100010000000001000000010000111100),
.INIT_2E(256'b0000000000001011000000000000010100000000000011110000000000000101000000000000111100000000000011110000000000001111000000000000101100000000000010010000000000001101000000000000100101000000000010100000000000000010010000000000100011000000000000011000000000001000),
.INIT_2F(256'b0101101000111111101111000011111101111110000111101111111100001100010111111100000011111111000000001111111010100010011111110100000011111110100100010111110100111001101111100010001101001100010001100011100000100010000111000111101000000011100001001000111000000011),
.INIT_30(256'b1111111111111100111111111111110000011111111111000000000111111100000000001111110000110000011111000001100001111100000100000111110000010000011111000011000001111100101100000111110000010000011111000000100001111100000100000111111000100000111111100000000111111111),
.INIT_31(256'b0111000110001100101000111000100001000111100010000000111100010000000111100000000000111000000000000000000001001010000000010101010000000101111010000110000101110100000001101111100010001101111101000010011111101000101011111111010011111111111010001111111111110000),
.INIT_32(256'b1111100000000001011111100000000000101111100001010001111111100000001011111100000100010111111111001010111111110010000101011111110110101111111111100101010111111110101011111111111100111111111111110000111111111101000001111111111000000111111111010000000011111110),
.INIT_33(256'b0000010000000000000000010000000000000000011010000000000000000000000000000000000010000000000000000101000000000000000110110011000000000000001111110000000000000000100000000000000000000000000000001010000000000000010000000000000010100000000010101111111101011000),
.INIT_34(256'b0000100000000110001000000000110100000000000101100000000000001010100000000001000001000000001000000011000010100000000100000000000000000101000011000000101111111010000001011111010100101010111111101000010111111110101111111111010000101111110101110000000000001111),
.INIT_35(256'b1000000000000000010100000000000010000000000000000100000000000000100000000000000000111000000000000100101100000000101111100101000001111111100001101111111101000001111110101000011011111111000011101111100000001111100000110001101000000000011000110000000001000010),
.INIT_36(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111110000000000000001000000000000000011101100000000001111111100010000),
.INIT_37(256'b1111111010101000111111111111000011111111101010101111101111010000111110011110101011111111111101001111111100111010111101010010110111111110101101101111010100001001111111101000010111110101000000100011111000000000111111010000000011100110100000001111010100000000),
.INIT_38(256'b1111100011100000111100000100000011100010101010001100011111000000100011111010100000011111110000000000111110010000010111110100000000111110100000000111111100000000111110101000001011111111000000101111101010000101111111010100111011111110101011101111111101111100),
.INIT_39(256'b0000011011111010000110111111010001000111111110001000111111110100001111111110100011111111111100101111111111101000111111111111000001011111101010001111111111110000010111111110000111111111001101011111101001111110110100111111111110000111111110100011111111111111),
.INIT_3A(256'b0000010101111011000000001011111100000000011111111000000010101111100000000111111100100000101011110001000001011111000000000011111111000010000111111110001000101111111100011001111111111000001011111111110000110111111111100000101111111111100001111111111111000001),
.INIT_3B(256'b0101110001111000100111100011000100111110001100011011111000100001001111000010000100111100000001010111111100000011011111100000001101111111100001111111111100000011111111111000001111111111111000111111111111000011111111111110101111111111111101111111111111111011),
.INIT_3C(256'b1110001001010101110000000010001011000100010001111000100000100011000000000100011000010000001010100010000001010000000000010100001101000101000111111001010001111111010100011111111111000111111111111000101111111111000101111111111100001011111111110001011111111111),
.INIT_3D(256'b0000000000000000000100000000000010001000000000001000110000000000110000000000000011100010000000001111000000000000111100010000000011111000110000001111110001100000111111100011000011111111000110001111111110001100111111111100011011111111111000111111111111110001),
.INIT_3E(256'b1111000010000000111000110000000011100000000000001100000000000000100011000000000010001000000000000001100000000000000100000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000001000000000000000100000000000000),
.INIT_3F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram4 (
      .DIA(dia[4]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4]),
      .SSRA(ssra),

      .DIB(dib[4]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(256'b1100000000000000110000000000000011000000000000001100000000000000110000000000000111000000000000011100000000000000110000000000000011000000000000011000000000000011100000000000000110000000000000011000000000000111000000000000001100000000000001110000000000000111),
.INIT_01(256'b1000011111111111010000111111111100100001111111110000000111111111000000001111111100000000011111110000000101111111000000001111111100000000001111110000000001111111000000000001111100000000010111110000000000001111000000000000111100000000000001110000000000011111),
.INIT_02(256'b1110100000000000101101000000000001101000000000001101000000000000111010100000000001010000000000001110101000000101010100000000111110101000000011110100000000011111101010001111111101000000111111111000011111111111010101111111111111011111111111110111111111111111),
.INIT_03(256'b1111111110111111111111111011111111111111101111111111111110111111111111110111111111111111011111111111111101111111111111111111111111111110111111111111111111111111111111010111111111111110001111101111100000010101111101000000101011110000000000011110100000000010),
.INIT_04(256'b1111110000010000111110101000010011111111010000101111101010000011111111110100000111111110100000001111111101000000111111101010000011111101000000001110101010100000110101010000000010110000101000001100000000000000111110000000000011111000000000001111111100000000),
.INIT_05(256'b1111111111011111101111100111111101110011111111110011111111111111111111111111110111111111111111111111111111111101111111111111111111111111111111011111111111111111111111111111110111111111111101011111111110010111111111001011111110001001111111110111111111111111),
.INIT_06(256'b0111111111111111111111111110111111111111111101111111111111110111111111111111111111111111111111111111111111110111111111111111111111111111101111111111111010111111111100101111111110010111111111110111111111111111111111111111111111111111111111111111111111111110),
.INIT_07(256'b1111111111111111111111111111111100011001111111111111111110111111111111111001011111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_08(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111000001111111111111100000111111111111110000),
.INIT_09(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111100011111111110000011111110000000111110000101010111111),
.INIT_0A(256'b1111111111111111111111111111111111111111111111011111111111110011111111111111000111111111111100001111111111111000111111111110100011111111100011001111110011110100000111111111110011111111111110101111111111111110111111111111110111111111111111111111111111111110),
.INIT_0B(256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111011111111111100010111110001111100000010001111110010000011111111001101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0C(256'b1010000010101000100000000010000010000000000110100000000101111110000000001011111100000101011111110000000010101111000001011111111110000000101011110010000101111111110010001010111111110010111111111111110010111111111111110111111111111111110101111111111111111010),
.INIT_0D(256'b0000000010111111000000000010111100000000000110010000000010101111000000000101111100000010101111110000000001010111100000001011111101000000010101111000000000111111111110000001111111110110000011111111110101000101111111111010111111111111111100111111111111111111),
.INIT_0E(256'b1111111110100111111111101111111111111101111111111111101111111111111100111111111111110011111111111110010111111111110010110111111100000101111111110000001010111111000101011111111100000010111100010001010111100011000000101101111100000001001111110000001000111111),
.INIT_0F(256'b0000000001111111000000000011111000000000011111010000001011111111000000111111111100000001111111110000101110111111000001111111111101011110111111111001111011111111001111110111111101111111111111011111111111011010111111111110100011111111111110001111111111111111),
.INIT_10(256'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000001000000000000000010000000000000000000000000000000110110000000000010111000000000001100100000000001111),
.INIT_11(256'b1111111111111111111111111111111111111111111111111111111111111110111111111111110111111111111110111111111111110111111111111110111111111111110111111111111111011111111111111011111101111111011101111101111111111111111011100101011111110110001011111111110000010111),
.INIT_12(256'b1111111100010111101011110010111111111111110111111010111111011111010101111000111110101111111011110001010101011110001010111100111010000101010111111010101011000111000000010100110011000010100000100000000001000101000000001000000001000000010000000010000000000000),
.INIT_13(256'b1111111101000001111111111000000011111111010000101111111101000010111111110110001111111111101111101111111110110010111111111111100011111111111110100111111111011000001111111101110001111111110111111101111111011110101111111111111011011111111111101111111110001110),
.INIT_14(256'b1111110111111110111111011111111011111111111111001111110111111101111110011111110011111111111111011111101111111100111111111111110111110011111111011111011111111111111111111111111011111111111111111111111111111111110111111111111110011111111111111111111111111111),
.INIT_15(256'b1111100111111111111111011111111111111101111111111111110011111111111111011111111111111110111111111111111011111111111111000111111111111100111111111111110001111111111111000011111111111101111111111111110100111111111111101001111111111110111111111111111011011111),
.INIT_16(256'b1011110011111111111111010111111101111110011111111111111101111111011111111011111111111110111111110111111001111111111111110011111111111111100111111111111110011111111111110111111111111111011111111111111111011111111111111101111111111111111010111111111111111011),
.INIT_17(256'b0111010100001111000111110000111111101011101111111111111110101111111110001001111111111110100011111111110011011111111111111101111111111111110111111111111100001111111111111100111110111111100011111111111111111111101111111101111111111111111111111011111111111111),
.INIT_18(256'b1000000000000101100000000000001011000000000001011100000000000000000000000000010100000000000000111000000000000010110000000000001111000000000001011100000000000011100000000000101111100000000001111100000000010111111100000010111111111000010111111110101110111111),
.INIT_19(256'b0000000001100101000000001100100100000000010000110000000001000011000000001100001100000000100010100000000010011101000000000101101000000000010100010000000000000010000000000101000100000000010100100000000000110001000000000010001000000000000000010000000000100010),
.INIT_1A(256'b0000000000000010000000000000101000000000000011100000000000011111000000000001111100000000001011110000000000011111000000000001111100000000111111110000000001111111000000000111111100000010111111110000010111111111000100111111111101011111111111111101111111111111),
.INIT_1B(256'b0000000000000000000000000001100000000000000010001000000000000110000000000000011001100000000000101010000000000010110100000000001001110100000000001011000000000000011110100000000000111100000000000001111000000000000011100000000000000110000000000010011000000000),
.INIT_1C(256'b1100000000011001110000000000000011010000000000001100000000000000111100000000000011101000000000001110000000000000111110000000000011110000000000001111110000000000111110100000000011111100000000001111111100000000111111111110000011111111101111111111111111110000),
.INIT_1D(256'b0000000000000000000000000000011100000000000000110000000000000010000000000000000101000000000000100000000000000000010000000000000010000000000000110000000000000010000000000000010000000000000000000000000000001000000000000001000000000000000010000000000000010100),
.INIT_1E(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111),
.INIT_1F(256'b1000000001101111100000000000111110000000010011110000000000001111000000000100111110000000010011110000000000101111000000000000111110000000001011111000000000001111100000000010111110000000001011111000000000011111100000000000011110000000000101111000000000000111),
.INIT_20(256'b1111001100100000110101111100000010100011100000001100001100000110000010110001100010011011000000001110001100100000010000011000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100),
.INIT_21(256'b1101000000000011110000000000001010000000000000010010000000000001100000000000011110000000000000011000000000000011000000000000111100000000000011101000000000010110100000000001011000000000000111110100000000111111100110011101111111010001001111101111000011111110),
.INIT_22(256'b1010000000000011110000000000000111010000000000001111000000000000111100000000000011101000000000001111000000000000111110000000000011111000000000001111000000000000111100000000000011110000000000001111010000000000111101000000000011110100000000001111010000000000),
.INIT_23(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111100001011111111110110001011111111),
.INIT_24(256'b0000000011111111000010111111111100001011111111110000101111111111000010001111111100001000111111110000100111111111000010011111111100000001111111110000000111111111000000010111111100000000011111110000100001111111000011001111111100000100101111110000000000111111),
.INIT_25(256'b1111111111111111111111111111111111111111111110101111111111101000111111111101000011111111100101111111111010100000111111101000000011111010000000001110100000000000110000000000000010100000000000001100000000000000110000000000000000000000000000001000000000000000),
.INIT_26(256'b1111111100100000111111110011000011111111001100001111111100110000111111110101000011111111011100001111111010110000111111110111000011111110111100001111100011110000111101111111000010001101111100001111111111110000001111011111000000000010111100001101110101110000),
.INIT_27(256'b1000001000001111011110011000111111111100000011111111111010011111111111101001111111111110100111111111111010011111111111101001111111111110100111111111111010011111111111101001111111111110100111111111111010011111111111100001110111111110000111011111111000001100),
.INIT_28(256'b1111110000101111111111001110111111110000010011111111100111111111111000101101111111100101111111111100100110011111100101111001111100111111110111111111111111111111111111111111111111111111110011111111111111101111111111111110011111111111111100111111111111111100),
.INIT_29(256'b1111111111111011111111111011101111111111101111111111111101111101111111111111110111111111011111111111111101110111111111101111011111111110111101011111111111111001111111011110100111111101111010011111110111111011111110111101100111111111110111111111111111010011),
.INIT_2A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111011111111011100011111111011100000001111111110000001011111100000000011111000110100001111111101010000001111111000000010110),
.INIT_2B(256'b1111111111111111011111111110011101111111111101110111111111111011001111111111011110111111111110111111111111111011101111111111111111011111111111111101111111111111111111111111111111001111111111111111111111111111110111111111111101100111111111111111111111111111),
.INIT_2C(256'b1000000101111101100000000111111010000000111111010000000010111111110000101011001111000001111011111110001011000111011100010100111101100010111001110011000111101111011110101110001100110001111111110101101111110011101011111111011101011001111110011011110111111001),
.INIT_2D(256'b1000000000001000100000000000100010000000000010001000000000001000100000000000100010000000000010001000000000001001100000000000100111000000000000101100000000001100100000000000011111000000000000001010000000000000111000000000001011111000000001111111010000010011),
.INIT_2E(256'b0000000000001011000000000000010100000000000011110000000000000101000000000000111100000000000011110000000000001011000000000000111100000000000010010000000000001011000000000000110100000000000011000100000000000101010000000000111001000000000001101000000000001111),
.INIT_2F(256'b1111100111111111111111011111111111111110111111111111111101111111111111111011111111111111001111111111111010011100111111110101101101111110100001101011110100011110010111100011110000111100011110000001100010111000000001011111110000001100100001100000001000000010),
.INIT_30(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111011111111111111101111111111111110111111111111101011111111111001001111111111111100111111111111111011111111111111011111111111111011111111111110111111111111111),
.INIT_31(256'b0110111111110000000111111111100000111111111100001111111111101000111111111111000011111111110100001111111110000000111111100000000011111001000000001000000010000000000001010000000010001010000000000011000000000000110100000000000001000000000000000000000000000000),
.INIT_32(256'b0001011111111111100001011111111111010001011111111110000001011111110100000010111111101000000010110101000000001101111010100000001001010000000000011010101000000001010100000000000001000000000000001101000000000000111100000000000011111010000000001111111000000000),
.INIT_33(256'b1111110111111111111111110111111111111111111001111111111111111111111111111111111101111111111111111100111111111111111001110000111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111100110111),
.INIT_34(256'b1001011111111000110111111111001111111111111010011111111111110001111111111110001111111111110001111101111110011111111101111111111111111100111100001111111111111010111111111111010111111111111111101111111111111111011111111111100111100000000110001111111111110000),
.INIT_35(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111001111111001111101111111111110111111111111111110111111111111100111111111111100011111111111110000000000001110000111111111111000001111111110010001),
.INIT_36(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111100001111),
.INIT_37(256'b1011111111111111110111111111111111101111111111111111001111111111111111011111111111111110111111111111111110111111111111111100111111111111111110111111111111111001111111111111110011111111111111100111111111111111110111111111111111101111111111111111001111111111),
.INIT_38(256'b1111111100111111111111100111111111111110111111111111111111111111111111111111111111111111111111111100111111111111100111111111111111111111111111110111111111111111011111111111111111111111111110101111111111110101111111111110111011111111111111111111111111011101),
.INIT_39(256'b1111100011111111111000111111111110000111111111110000111111111111001111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111010111111111111011111111110001101111110001111111111000111111111100000111111111110011111111111111),
.INIT_3A(256'b0000010101111001000000001011111000000000011111110000000010101111010000000111111111100000101011111111000001011111111100000011111111111000000111111111110100101111111111101001111111111111100011111111111111000111111111111111101111111111111110011111111111111111),
.INIT_3B(256'b0101111111111111000111011111111110111101111111101011110111111101001111011111111100111101111110010111111011111011011111101111111101111111011110111111111101111011111111111011101111111111110110111111111111011011111111111110001111111111111100111111111111111111),
.INIT_3C(256'b1111110001010101111111000010001011111000010001111111000000100011111100000100011111100000001011001100000001100000110000011000001110000110000111110001100001111111011000011111111110000111111111110000101111111111000101111111111100001011111111110001011111111111),
.INIT_3D(256'b1111000000000000111000000000000011111000000000001111000000000000111110000000000011111110000000001111111100000000111111101000000011111111000000001111111110000000111111111100000011111111111000001111111111110000111111111111100011111111111111001111111111111110),
.INIT_3E(256'b1111111000000000111111000000000011111110000000001111100000000000111100000000000011111000000000001110000000000000111100000000000011100000000000001100000000000000111000000000000011000000000000001000000000000000110000000000000010000000000000001000000000000000),
.INIT_3F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram5 (
      .DIA(dia[5]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[5]),
      .SSRA(ssra),

      .DIB(dib[5]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[5]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000010000000000000001000000000000001100000000000000110000000000000011000000000000011100000000000001110000000000001111),
.INIT_01(256'b1011111111111111010111111111111100101111111111110000011111111111000000111111111100000001111111110000000011111111000000000111111100000000011111110000000000111111000000000011111100000000010111110000000000011111000000000000111100000000000011110000000000010111),
.INIT_02(256'b0000100000000000001101000000000001101000000000001101000000000000111010100000000001010000000000011110101000000011010100000000011110101000000111110100000000111111101010000111111101000001111111111000001111111111010011111111111110111111111111111111111111111111),
.INIT_03(256'b1111111111000000111111111100000011111111110000001111111111000000111111111000000011111111100000001111111110000000111111110000000011111111000000001111111000000000111111101000000011111101110000011111111111101010111110111111010111111111111111101111011111111101),
.INIT_04(256'b1111110000001111111110101000001111111111010000011111101010000010111111110100000111111110100000001111111101000000111111101010000011111101000000001110101010100000110101010000000000110000101000001110000000000000111100000000000011111100000000001111111000000000),
.INIT_05(256'b0000000000011111010000000111111110000011111111110011111111111111111111111111110111111111111111111111111111111101111111111111111111111111111111011111111111111111111111111111110011111111111100111111111110001111111111000111111110000111111111111111111111111111),
.INIT_06(256'b0111111111101111111111111110011111111111111101111111111111110111111111111111111111111111111111111111111111110111111111111110111111111111100111111111111001111111111100011111111110001111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_07(256'b1111111111111111111111111111111111100001111111111111111000111111111111111110011111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_08(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111100000000011111110000000000001111),
.INIT_09(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111100011111111111000001111010101000000),
.INIT_0A(256'b1111111111111111111111111111111111111111111100111111111111110000111111111111000011111111111100001111111111110000111111111111000011111111111100001111111100001000111000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000001),
.INIT_0B(256'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011111111110011111111111111100011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0C(256'b0001111110010111011111111110111111111111111110011111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111011111111111111111011111111111111111011111111111111111011111111111111111001111111111111111100),
.INIT_0D(256'b1111111110000000111111111110000011111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111011111111111111111011111111111111111001111111111111111100111111111111111111001111111111111111),
.INIT_0E(256'b0000000000111111000000001111111100000001111111110000001111111111000001111111111100011111111111110011111111111111011111111111111101111111111111111111111111111111111111111111111011111111111110111111111111110111111111111110111111111111110111111111111110111111),
.INIT_0F(256'b1111111101111111111111111111111111111110111111101111111111111000111111011111000011111011111000001111111111000000111111110000000010101111000000000111111100000000111111111000000111111111100000001111111111100001111111111111011111111111111111011111111111111110),
.INIT_10(256'b1111111111111111011111111111111101111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111100111111111111110011101111111111011100111111111101110011111111110111),
.INIT_11(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111001111111111111000111111111111000011111111111000001111111111100000111111111100000011111111100010000011111100000000000111111010100000001111110100000000001111101000),
.INIT_12(256'b0000000011100000010100001010000000000000001000000101000001100000101010000101000001010000001100001110101010100000110101000010000001111010101100010101010100110001111111101011100110111101011110110111111110111110011111110111111101111111101111110001111111111111),
.INIT_13(256'b1111111110000000111111110000000011111111100000111111111110000010111111111000000011111111110001011111111111000001111111111100001111111111110000111111111111100001011111111110000110111111111000010111111111100000010111111110000000011111111000000011111111110000),
.INIT_14(256'b0000000111111100000000011111110000000001111111100000001111111110000001111111111000000111111111100000001111111110000000111111111000001111111111100000011111111110000001111111111100011111111111110000111111111111000111111111111100111111111111110111111111111111),
.INIT_15(256'b0000010000000000000000000000000000000000000000000000000100000000000000010000000000000010000000000000001000000000000000101000000000000010100000000000001000000000000000100100000000000010010000000000001000000000000000010010000000000001001000000000000100000000),
.INIT_16(256'b0011110100000000001111111000000011111110100000001111111010000000011111101100000001111111110000001111111101000000111111110000000011111111001000001111111100100000111111111010000011111111101000001111111110000000111111111111000011111111111111111111111111111111),
.INIT_17(256'b0111001000100000000001000010000000000100001000000000001000100000000000100000000000000000000000000000000100000000000000000000000000000000100000000000000010010000000000000101000000000000010100000000000000110000000000000011000000000000000100000000000000010000),
.INIT_18(256'b0100000000000000010000000000000001000000000000000100000000000001100000000000000110000000000000001000000000000001100000000000001110000000000000011000000000000111110000000000001111000000000011111110000000000111110000000000111111110000000111111111001101111111),
.INIT_19(256'b0000000000000000000000001000100000000000100010000000000010001000000000000000100000000000000000000000000000010000000000000101000000000000010100000000000001010000000000000000000000000000000000000000000000100000000000000010000000000000001000000000000000000000),
.INIT_1A(256'b1000000000000011000000000000011100000000000011110000000000000111000000000001111100000000000111110000000000011111000000000111111100000000001111110000000001111111000000001111111100000011111111110000011111111111000001111111111100101111111111111011111111111111),
.INIT_1B(256'b0000000000010100000000000000110000000000000001000000000000000000010000000000000000100000000000000000000000000000000010000000000010000000000000000100010000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000010000000000000),
.INIT_1C(256'b1111000000010001111100000001001011110000000000001110000000000000111000000000000011110000000000001111100000000000111100000000000011111100000000001111100000000000111111100000000011111111000000001111111010000000111111110100000011111111110100001111111111111111),
.INIT_1D(256'b0000000000000100000000000000001000000000000000110000000000000010000000000000001001100000000000010010000000000011010000000000001110000000000000100000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000011000),
.INIT_1E(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_1F(256'b0000000001111111000000000011111100000000011111111000000001111111100000000011111110000000001111110000000000011111000000000001111100000000001111110000000000111111000000000001111100000000000111110000000000001111000000000000111100000000000111110000000000011111),
.INIT_20(256'b1111111111000000111000000000000011000000000000001000000000000100100010000000000000010100000000000100000000000000000000001000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_21(256'b1110000000000000110000000000000111100000000000111000000000000001010000000000000110000000000001110000000000000011000000000000001100000000000011110000000000000111000000000001111100000000001011101100000001011110110000001011111011100000111111111111111111111111),
.INIT_22(256'b1100000000000000110000000000000011100000000000001111000000000000111000000000000011110000000000001111100000000000111110000000000011110000000000001111100000000000111110000000000011111000000000001111100000000000111110000000000011111000000000001111100000000000),
.INIT_23(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111110110000111111111),
.INIT_24(256'b0000100111111111000010011111111100001001111111110000100111111111000010011111111100001001111111110000100011111111000010001111111100001000111111110000100011111111000010001111111100001000111111110000000011111111000001000111111100000100011111110000010001111111),
.INIT_25(256'b1111111111111111111111111111111111111111111111001111111111110000111111111110000011111111110110001111111101000000111111010000000011111000000000001111100000000000111100000000000011100000000000001100000000000000000000000000000010000000000000000000000000000000),
.INIT_26(256'b0000000000010000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000101100000000000011110000000000000111000000000001111100000000000011110000001111011111000001111111111100000110000111110000000000001111000000011110011100000),
.INIT_27(256'b0000000100001111000000001000111100000000100011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011100000000000001111000000001000111000000000100011000000000010011110),
.INIT_28(256'b0000010001111000000001000110000000001000111100000000100011000000000100011100000000010011111000000010011111100000010011111110000001111111111000001111111111100000111111111100000011111111111100001111111111100000111111111111000011111111111110001111111111111110),
.INIT_29(256'b0000000001000000000000000000000000000000000000000000000010000010000000001000001000000000000000100000000000001010000000010000101000000000000010000000000000001100000000100001110000000000000111000000000000011110000001000011111000000100001110000000010000111000),
.INIT_2A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111100000000111111100000000011111100000000000111110000000000001111111110100000111100000110000011110000001000001111),
.INIT_2B(256'b0000000000010000100000000001000010000000000000000000000000001000010000000000110001000000000001000100000000000100000000000000000000100000000000000000000000000000000000000000000000110000000000000011000000000000001000000000000000111000000000000011100000000000),
.INIT_2C(256'b1000000011111110100000001111110000000000011110100100000001110100000000000111010000100000001110000000000000111000100100000011100010010000000100001100000000010000100010000001110011001000000011001010000000001000010101000000100010100100000001100100000000000110),
.INIT_2D(256'b1111111111111000111111111111100011111111111110001111111111111000111111111111100011111111111110001111111111111000111111111111100011111111111110001111111111110000101111111111101110111111111111001111111111111110110111111111111011101111111111011111111111110111),
.INIT_2E(256'b1111111111110100111111111111101011111111111100001111111111111010111111111111000011111111111100001111111111110100111111111111010011111111111100101111111111110010111111111111000011111111111100011111111111111001111111111111000011111111111110001011111111110000),
.INIT_2F(256'b0000011111111111000000111111111100000001111111110000000011111111000000000111111100000000111111110000000101111111000000001011110000000001011110001000001011100000110000011100000011100011100000001111011100111000111100101000000111111001011110001111101111111100),
.INIT_30(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111110000111111111111000011111111111100001111111111110000111111111111110011111111111111111111111111111111111111111111111011111111111111011111111111110011111111111111),
.INIT_31(256'b0001111111111111011111111111011111111111111101111111111111111111111111111110111111111111111111111111111111011111111111111011111111111110011111111111111011111111111110011111111101110011111111111100011111111111000111111111111101111111111111111111111111111111),
.INIT_32(256'b1111000000000000111111000000000011111111000000001111111111000000111111111110000011111111111110001111111111111100111111111111111011111111111111111111111111111111111111111111111101111111111111110001111111111111000001111111111100000011111111110000000011111111),
.INIT_33(256'b0000001111111111000000001111111100000000000111110000000000000000000000000000000000000000000000001100000000000000111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100001111),
.INIT_34(256'b1100011111111110111111111111111011111111111111011111111111111011111111111111011101111111111011110001111110111111000011111111111100000011111111110000000000000101000000000000101000000000000000010000000000000000000000000000000111100000000111111111111111111111),
.INIT_35(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111110000000001111110000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000001111111111101000),
.INIT_36(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111),
.INIT_37(256'b0011111111111111000111111111111100001111111111110000001111111111000000011111111100000000111111110000000000111111000000000000111100000000000000110000000000000110000000000000001100000000000000010000000000000000110000000000000011100000000000001111000000000000),
.INIT_38(256'b1111111110111111111111110111111111111100111111111111101111111111111101111111111111101111111111111110111111111111110111111111111110111111111111111111111111111111011111111111111011111111111110011111111111110010111111111110000111111111111000011111111111000011),
.INIT_39(256'b1111111100000000111111000000000011111000000000001111000000000000110000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000101000000000000000000000000001110000000001111111000000111111111100000111111111110011111111111111),
.INIT_3A(256'b0000010101111000000000001011111000000000011111110000000010101111100000000111111111000000101011111110000001011111111110000011111111111100000111111111111000101111111111110001111111111111110011111111111111100111111111111111001111111111111111011111111111111110),
.INIT_3B(256'b0010001111111111011000111111111001000011111111100100001111111111110000111111110111000011111111011000000111111111100000011111101110000000111110110000000011111011000000000111101100000000001110110000000000111011000000000001101100000000000010110000000000000011),
.INIT_3C(256'b1111111110101010111111111101110111111111101110001111111111011100111111111011100011111111110100001111111110000000111111100000001111111000000111111110000001111111100000011111111100000111111111110000101111111111000101111111111100001011111111110001011111111111),
.INIT_3D(256'b1110000000000000111100000000000011110000000000001111100000000000111111000000000011111100000000001111111000000000111111110000000011111111100000001111111111000000111111111110000011111111111100001111111111111000111111111111110011111111111111101111111111111111),
.INIT_3E(256'b1111111100000000111111100000000011111100000000001111110000000000111110000000000011110000000000001111000000000000111000000000000011100000000000001110000000000000110000000000000011000000000000001100000000000000100000000000000010000000000000001000000000000000),
.INIT_3F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram6 (
      .DIA(dia[6]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[6]),
      .SSRA(ssra),

      .DIB(dib[6]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[6]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_01(256'b0111111111111111101111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111101111),
.INIT_02(256'b1111011111111111110010111111111110010111111111110010111111111111000101011111111110101111111111110001010111111111101011111111111101010111111111111011111111111111010101111111111110111111111111110111111111111111101111111111111101111111111111111111111111111111),
.INIT_03(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_04(256'b0000001111111111000001010111111100000000101111110000010101111101000000001011111000000001011111110000000010111111000000010101111100000010111111110001010101011111001010101111111111001111010111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_05(256'b1111111111100000111111111000000011111100000000001100000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001100000000000011110000000001111111000000111111111101111111111111111111111111111111),
.INIT_06(256'b1000000000011111000000000001111100000000000011110000000000001111000000000000011100000000000001110000000000001111000000000001111100000000011111110000000111111111000011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_07(256'b0000000000000000000000000000000011111110000000001111111111000000111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_08(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_09(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_0B(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111100000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_0C(256'b1100000001111111100000000001111100000000000001110000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000111100000000000011111100000000001111111100000000111111111100000011111111111110001111111111111111),
.INIT_0D(256'b0000000001111111000000000001111100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001110000000000000111100000000000011111100000000001111111110000000111111111111000011111111111111111111111111111111),
.INIT_0E(256'b1111111111000000111111110000000011111110000000001111110000000000111110000000000011100000000000001100000000000000100000000000000010000000000000000000000000000000000000000000000100000000000001110000000000001111000000000001111100000000001111110000000001111111),
.INIT_0F(256'b0000000011111111000000001111111100000001111111110000000111111111000000111111111100000111111111110000011111111111000011111111111100011111111111110011111111111111011111111111111011111111111111101111111111111100111111111111100011111111111111101111111111111111),
.INIT_10(256'b0000000000000000100000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011000000000000001100000000000000111010000000000011111000000000001111),
.INIT_11(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_12(256'b0000000000001111000000000101111100000000011111110000000000111111000000000011111100000000000111110000000000011111000000000001111100000000000011100000000000001110000000000000011000000000000001001000000000000000100000000000000010000000000000001100000000000000),
.INIT_13(256'b1111111111111111111111111111111111111111111111001111111111111100111111111111110011111111111110001111111111111100111111111111110011111111111111001111111111111110111111111111111001111111111111100011111111111111001111111111111100111111111111110001111111111111),
.INIT_14(256'b0000001111111111000000111111111100000011111111110000001111111111000000111111111100000011111111110000011111111111000001111111111100000111111111110000111111111111000011111111111100001111111111110001111111111111001111111111111101111111111111111111111111111111),
.INIT_15(256'b0000001000000000000000100000000000000010000000000000001000000000000000100000000000000001000000000000000100000000000000010000000000000001000000000000000110000000000000011000000000000001100000000000000111000000000000011100000000000001110000000000000111100000),
.INIT_16(256'b0111111000000000011111100000000001111111000000000111111100000000111111110000000011111111000000001111111110000000111111111100000011111111110000001111111111000000111111111100000011111111110000001111111111100000111111111110000011111111111100001111111111111111),
.INIT_17(256'b1000111111000000000000111100000000000011110000000000000111000000000000011110000000000001111000000000000011100000000000001110000000000000011000000000000001100000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_18(256'b1000000000000000100000000000000010000000000000001000000000000000110000000000000011000000000000011100000000000001110000000000000111000000000000111100000000000011110000000000011111000000000001111100000000001111111000000001111111100000001111111111110011111111),
.INIT_19(256'b0000000011111000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1A(256'b0000000000000111000000000000011100000000000001110000000000001111000000000000111100000000000111110000000000111111000000000011111100000000011111110000000011111111000000011111111100000001111111110000001111111111000011111111111100011111111111110111111111111111),
.INIT_1B(256'b0000000000001000000000000000000000000000000000000000000000000000100000000000000011000000000000001111000000000000111100000000000011111000000000001111100000000000111111000000000011111100000000001111110000000000111111000000000011111100000000001101110000000000),
.INIT_1C(256'b1110000000001110111000000000110011100000000000001111000000000000111100000000000011110000000000001111000000000000111110000000000011111000000000001111110000000000111111000000000011111110000000001111111100000000111111111000000011111111111000001111111111111111),
.INIT_1D(256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000110000000000000011100000000000001100000000000000100000000000000010000000000000001000000000000001100000000000000110000000000000111000000000000111100000000000111110000000000100000),
.INIT_1E(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_1F(256'b0000000000111111000000000111111100000000001111110000000000111111000000000011111100000000001111111000000000111111100000000011111110000000000111111000000000011111100000000001111110000000000111111000000000011111100000000001111110000000000011111000000000001111),
.INIT_20(256'b1111111111111111111111111111111111111111111111111111111111111000111101111111000011100011111000001000001111000000100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011),
.INIT_21(256'b1110000000000001111000000000000111000000000000011100000000000011100000000000001100000000000000110000000000000111000000000000011100000000000001110000000000001111000000000000111110000000000111111000000000111111111000000111111111111111111111111111111111111111),
.INIT_22(256'b1100000000000000111000000000000011100000000000001110000000000000111100000000000011110000000000001111000000000000111100000000000011111000000000001111100000000000111110000000000011111000000000001111100000000000111110000000000011111000000000001111100000000000),
.INIT_23(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111),
.INIT_24(256'b0000011111111111000001111111111100000111111111110000011111111111000001111111111100000111111111110000011111111111000001111111111100000111111111110000011111111111000001111111111100000111111111110000011111111111000000111111111100000011111111110000001111111111),
.INIT_25(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111110000000111111100000000011111100000000001111000000000000111000000000000011000000000000001000000000000000100000000000000000000000000000000000000000000000),
.INIT_26(256'b0000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000001111000000000000111100000000000111110000000000111111000001111111111100000111111111110000011111111111000000000001111100000),
.INIT_27(256'b0000000011111111000000000111111100000000011111110000000001111111000000000111111100000000011111110000000001111111000000000111111100000000011111110000000001111111000000000111111100000000011111110000000001111110000000000111111000000000011111100000000001111100),
.INIT_28(256'b0000001111110000000000111111000000000111111000000000011111100000000011111110000000001111110000000001111111000000001111111100000011111111110000001111111111000000111111111110000011111111111000001111111111110000111111111111100011111111111111001111111111111111),
.INIT_29(256'b0000000000111100000000000111110000000000011111000000000001111100000000000111110000000000111111000000000011111100000000001111110000000001111111100000000111111110000000011111111000000011111111100000001111111100000000111111110000000011111111000000001111111100),
.INIT_2A(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001011111111100000001111111110000000111111111),
.INIT_2B(256'b0000000000001100000000000000110000000000000011001000000000000100100000000000000010000000000000001000000000000000110000000000000011000000000000001110000000000000111000000000000011100000000000001110000000000000111100000000000011110000000000001111000000000000),
.INIT_2C(256'b0111111111111111011111111111111101111111111111000011111111111000001111111111100000011111111100000001111111110000000011111111000000001111111110000000111111111000000001111111100000000111111110000000011111111100000000111111110000000011111111000000001111111100),
.INIT_2D(256'b1000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111110000000000000011000000000000011100000000000001111000000000000111110000000000111111100000001111),
.INIT_2E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000011000000000000001100000000000000110000000000000011100000000000001110100000000000111),
.INIT_2F(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111001111111111111100011111111111110000111111000111000011110000000000000110000000000000010000000000),
.INIT_30(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111100001111111111110000111111111111000111111111111100111111111111111111111111111111),
.INIT_31(256'b1111111111111000111111111111100011111111111110001111111111110000111111111111000011111111111000001111111111100000111111111100000011111111100000001111111100000000111111100000000011111100000000001111100000000000111000000000000010000000000000000000000000000000),
.INIT_32(256'b0000111111111111000000111111111100000000111111110000000000111111000000000001111100000000000001110000000000000011000000000000000100000000000000000000000000000000000000000000000010000000000000001110000000000000111110000000000011111100000000001111111100000000),
.INIT_33(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111111),
.INIT_34(256'b0011100000000001000000000000000100000000000000110000000000000111000000000000111110000000000111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111000000000000000000000),
.INIT_35(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111111110000011111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111110000000000000111),
.INIT_36(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_37(256'b1100000000000000111000000000000011110000000000001111110000000000111111100000000011111111000000001111111111000000111111111111000011111111111111001111111111111111111111111111111111111111111111111111111111111111001111111111111100011111111111110000111111111111),
.INIT_38(256'b1111111111000000111111111000000011111111000000001111110000000000111110000000000011110000000000001111000000000000111000000000000011000000000000001000000000000000100000000000000100000000000001110000000000001111000000000001111100000000000111110000000000111111),
.INIT_39(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111110000000111111000000000011111000000000001100000000000000),
.INIT_3A(256'b1111101010000111111111110100000111111111100000001111111101010000111111111000000011111111010100001111111110100000111111111100000011111111111000001111111111010000111111111110000011111111111100001111111111111000111111111111110011111111111111101111111111111111),
.INIT_3B(256'b1111111111111111111111111111111111111111111111111111111111111110111111111111111011111111111111101111111111111100111111111111110011111111111111001111111111111100111111111111110011111111111111001111111111111100111111111111110011111111111111001111111111111100),
.INIT_3C(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111000001111111110000000111111100000000011111000000000001111010000000000111010000000000011110100000000001110100000000000),
.INIT_3D(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_3E(256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
.INIT_3F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)
    ) ram7 (
      .DIA(dia[7]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[7]),
      .SSRA(ssra),

      .DIB(dib[7]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[7]),
      .SSRB(ssrb)
      );
`endif 

endmodule //SPRIMG


module RAM_PICTURE (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [12:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [12:0] addrb
    );

`ifdef GENERIC_RAM
	srambDrsws #(
		.DATA_WIDTH(8),
		.ADDR_WIDTH(13)
	) ram (
		.DIA(dia),
      .WEA(wea),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa),

      .DIB(dib),
      .WEB(web),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob),
	);
	
`elsif ALTERA
	RAMB32_S8_S8 ram(
	   .DIA(dia),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa),
      .SSRA(ssra),

      .DIB(dib),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob),
      .SSRB(ssrb)
	);
`else
    RAMB16_S4_S4 #(
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0C(256'h00000000000000000000BA900000000000008760000000000000005432100000),
.INIT_0D(256'h0000000000000000003211100FEDC0BA098760005403201000F0E0D0000C0000),
.INIT_0E(256'h00000000000000000000000000000000000000000000007654D0000000000D00),
.INIT_0F(256'h0000000000000000800000000000000000000000000000000000000000000000),
.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_11(256'h00000000000000A0000000000000000000000000000000000000000000000009),
.INIT_12(256'h00000000000000C000000000000000000000000000000000000000000000000B),
.INIT_13(256'h00000000000000E000000000000000000000000000000000000000000000000D),
.INIT_14(256'h000000000000000000000000000000000000000000000000000000000000000F),
.INIT_15(256'h0000000000000000000000000000000000200000000000000000000000000001),
.INIT_16(256'h0000000000000000000000000000000000300000000000000000000000000000),
.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_19(256'h0000000000000000000000050000000000000000000000000000004000000000),
.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000098760),
.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000FEDCBA),
.INIT_22(256'h0000000000000009807600000000000000000000000000000000000000543210),
.INIT_23(256'h0000000000000002101000000000000000000000000000000000000000FEDCBA),
.INIT_24(256'h000000000000000CBA9000000000000000000000000000000000000000876543),
.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000210FED),
.INIT_26(256'h00000000000000E414056FC0C5B21C30925B1A0CEF309D0F4091484292090018),
.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_28(256'h000E8FAADD0E3EF93310025F905532500B3E2F3105C449C0DF2603B1F094879D),
.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2A(256'h00000000007E94457025F90EF055EFC5D04E10C51839D0F403EF941C54127EF3),
.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2C(256'h000000000000000000000000DF3E44F254417E7770D039EF2435C5044F254417),
.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2E(256'hEFA526E7726EFA9E5EC6EFA9E927EF6EFA52F8A9849BBA9210280B0BE1965213),
.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_30(256'h0000000000E9F20C56FC0E25650569704352058407E95202F603BE1840A9DD14),
.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_32(256'h010254F39F27F305840DF260CCC10F407E9D170F245204E107E9B31809001801),
.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_34(256'h000000000000000000000000000321C3E93415800BE1C07E17005665400B5D20),
.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_36(256'h000000000000000000000000000000000DF3E3B3F2E17154060DF3E3B3F29217),
.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_38(256'h0000E5EF057E1830F40541C0FF402565E0C569C01056180F40541C0FF402565E),
.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3A(256'h00000000000000000000000000000000004CF80CC533520F403BE1840C193503),
.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3C(256'h0000000000000000000000000000000000035B540B5254092045B3120435AF20),
.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3E(256'hDDDDDDDDDDDDDDDDDDDD011020DF3EFE9545D1709380DDDDDDDDDDDDDDDDDDDD),
.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram0 (
      .DIA(dia[4*0+3:4*0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*0+3:4*0]),
      .SSRA(ssra),

      .DIB(dib[4*0+3:4*0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*0+3:4*0]),
      .SSRB(ssrb)
      );

    RAMB16_S4_S4 #(
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0D(256'h0000000000000000008888880111101101111000110110100100000000000000),
.INIT_0E(256'h0000000000000000000000000000000000000000000000888800000000000100),
.INIT_0F(256'h0000000000000000800000000000000000000000000000000000000000000000),
.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_11(256'h0000000000000080000000000000000000000000000000000000000000000008),
.INIT_12(256'h0000000000000080000000000000000000000000000000000000000000000008),
.INIT_13(256'h0000000000000080000000000000000000000000000000000000000000000008),
.INIT_14(256'h0000000000000090000000000000000000000000000000000000000000000008),
.INIT_15(256'h0000000000000000000000000000000000900000000000000000000000000009),
.INIT_16(256'h0000000000000000000000000000000000900000000000000000000000000000),
.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_19(256'h0000000000000000000000090000000000000000000000000000009000000000),
.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000099990),
.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000999999),
.INIT_22(256'h000000000000000AA0AA00000000000000000000000000000000000000AAAAAA),
.INIT_23(256'h000000000000000BB0BB00000000000000000000000000000000000000AAAAAA),
.INIT_24(256'h000000000000000BBBB000000000000000000000000000000000000000BBBBBB),
.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000CCCBBB),
.INIT_26(256'h2222222222222226662676622667664277666522667276267276667766277764),
.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_28(256'h2226666622227666776727767267777523767666266776626676276662776664),
.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2A(256'h2222222222666666727767266266666642666266666642672766676677676664),
.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2C(256'h2222222222222222222222226662776767767277722266667766662776767765),
.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2E(256'h5455554555154545555154545555551545554454554413233332245266676765),
.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_30(256'h2222222222276522676422767626667277662667266666276627666652376665),
.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_32(256'h2227666476676426652667622666267266666426776526662666666427776422),
.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_34(256'h2222222222222222222222222227666667776664266667666642767664263444),
.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_36(256'h2222222222222222222222222222222226662766656666652226662766657664),
.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_38(256'h2222266626666662672676626672767642266662626766267267662667276764),
.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3A(256'h2222222222222222222222222222222222766426667775267276666726666675),
.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3C(256'h2222222222222222222222222222222222276674266764276266666627666675),
.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3E(256'h2222222222222222222223333266626667666642242222222222222222222222),
.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram1 (
      .DIA(dia[4*1+3:4*1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*1+3:4*1]),
      .SSRA(ssra),

      .DIB(dib[4*1+3:4*1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*1+3:4*1]),
      .SSRB(ssrb)
      );
`endif
endmodule


module RAM_CHR (
    input [1:0] dia,
`ifdef GENERIC_RAM
    output reg [1:0] doa,
`else
	 output [1:0] doa,
`endif
    input wea,
    input ena,
    input clka,
    input ssra,
    input [14:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [12:0] addrb
    );

	 
	 
`ifdef GENERIC_RAM
	
	// Note, we will only ever be writing to port B
	// port A requires a selection on the address
	
	wire [7:0] tWire;
	
	srambDrsws #(
		.DATA_WIDTH(8),
		.ADDR_WIDTH(13)
	) ram (
		.DIA(0),
      .WEA(0),
      .CLKA(clka),
      .ADDRA(addra[14:2]),
      .DOA(tWire),

      .DIB(dib),
      .WEB(web),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob)
	);
	
	always @(addra[1:0],tWire)
  begin
    casex (addra[1:0])
    2'b00: doa <= tWire[1:0];
	 2'b01: doa <= tWire[3:2];
	 2'b10: doa <= tWire[5:4];
	 2'b11: doa <= tWire[7:6];
 
    // default: mem_data_rd_reg <= 0;
    endcase
  end
  
`elsif ALTERA
	RAMB32_S2_S8 ram (
      .DIA(dia),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa),
      .SSRA(ssra),

      .DIB(dib),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob),
      .SSRB(ssrb)
      );
	
`else
    RAMB16_S1_S4 #(
      .INIT_00(256'h00FFFFFF0000000000FFF7100000000000300000000000000000000000000000),
.INIT_01(256'h00FFEFCF000000000070300000000000CF0E00000000000000FFFF0E00000000),
.INIT_02(256'h0F00000000000000FF00000000000000F1000000000000000800000000000000),
.INIT_03(256'hF3F00000000000008F0E08000000000000000000000000FF00000000F1701000),
.INIT_04(256'h0000EFEFCF8F00000000F07030000000CF030000000000000F0C000000000000),
.INIT_05(256'h0000000000EFCF0F00000000007E3E0C000000FFEFC300000000F03000000000),
.INIT_06(256'h00000000008F0F0C0000000000FFF7F300FFFFCF00000000007E1C0800000000),
.INIT_07(256'h00000000FFEF8F0E00000000FFF7F3F00070301000000000000F000000000000),
.INIT_08(256'h006363F763F763630000000000C6C6C600810081818181810000000000000000),
.INIT_09(256'h00000000000381C000B366D683C6C6830060660381C066060081E7B0E386F3C0),
.INIT_0A(256'h00008181E7818100000081E7C3E78100000381C0C0C0810300C08103030381C0),
.INIT_0B(256'h0000060381C06000008181000000000000000000E70000000381810000000000),
.INIT_0C(256'h00C36660C16066C300E70381C06066C300E781818181838100C36667E7E666C3),
.INIT_0D(256'h0003030381C060E700C36666C70603C100C3666060C706E700C0C0E7C6C3C1C0),
.INIT_0E(256'h038181008181000000818100818100000083C060E36666C300C36666C36666C3),
.INIT_0F(256'h0081008181C066C3000381C060C08103000000E700E7000000C08103060381C0),
.INIT_10(256'h00C36606060666C300C76666C76666C700666666E76666C300C306E6A6E666C3),
.INIT_11(256'h00C36666E60666C300060606C70606E700E70606C70606E70087C6666666C687),
.INIT_12(256'h0066C6870787C6660083C6C0C0C0C0E300E78181818181E700666666E7666666),
.INIT_13(256'h00C36666666666C3006666E6E7676666003636B6B6F7773600E7060606060606),
.INIT_14(256'h00C36660C30666C3006666C6C76666C70063C6A6666666C300060606C76666C7),
.INIT_15(256'h003677F7B6B636360081C3666666666600C366666666666600818181818181E7),
.INIT_16(256'h00C70606060606C700E7060381C060E700818181C3666666006666C381C36666),
.INIT_17(256'hFF00000000000000000000002466C38100E36060606060E3000060C081030600),
.INIT_18(256'h00C3660666C3000000C7666666C7060600E366E360C3000000E70303C70363C1),
.INIT_19(256'hC360E36666E3000000030303C70303C100C306E766C3000000E3666666E36060),
.INIT_1A(256'h0066C687C6660606078181818183008100C38181818300810066666666C70606),
.INIT_1B(256'h00C3666666C300000066666666C700000036B6B6F763000000C3818181818183),
.INIT_1C(256'h00C760C306E300000006060667C600007060E36666E300000606C76666C70000),
.INIT_1D(256'h0063F7B6B63600000081C3666666000000E366666666000000C1030303C70303),
.INIT_1E(256'h00C08181078181C000E70381C0E70000C360E366666600000066C381C3660000),
.INIT_1F(256'hFFFFFFFFFFFFFFFF000000000064B61300038181E08181030081818100818181),
.INIT_20(256'h0F0E0800000000000000000000000C00000000000000FFFF00000000F1F03000),
.INIT_21(256'h000000000000FFEF0000000000703010000000000008000000000000000000CF),
.INIT_22(256'hF0F0F070707070700C080808000000007030303030101000000000000E0C0800),
.INIT_23(256'h10303030707070700C0C0C0C0E0E0E0E70F0F0F0F0F0F0F00E0E0E0E0E0C0C0C),
.INIT_24(256'h000000000000000E8F0000000000000000000000000000100000000000080808),
.INIT_25(256'h0F8F8F8F8FCFFFFFF9FFFFFFFFFFFFFF00000030000000000000000000000800),
.INIT_26(256'h08080000000070F0FFFFFFEFCFCFEFFF9FFFFFFFFFFFFFFFF0F1F1F1F1F3FFFF),
.INIT_27(256'hFFFFFFF7F3F3F7FF1010000000000E0F00000000000010F0000000000000080F),
.INIT_28(256'hCFCFCF8F0F080000F3F3F3F1F01000000000000000000808080CEFEFFFFFFFFF),
.INIT_29(256'h0F0F0F0F0F0000001C0C0ECFEFFFFFFF1030F7F7FFFFFFFF0000000000001010),
.INIT_2A(256'hF7F7FFFFFFFFFFFFFFFFEF0F0C0808081E1C0030B1FFFFFF7838000C8DFFFFFF),
.INIT_2B(256'hFFFFF7F030101010EFEFFFFFFFFFFFFF0F8F8FCFCFEFEFEFF0F1F1F3F3F7F7F7),
.INIT_2C(256'hCFEFFFFFFFFFFFFF0F0F0F0F0F0F0F0E0F0F0F0F0F0F0F0FFFFFFFFFFFFFFC3C),
.INIT_2D(256'h00000010101010008F8F8F0F0F0F0E0EF1F1F1F0F0F070700000000808080800),
.INIT_2E(256'hFFFF8D0C00B878F0000083838300000000000F0F0F0F0F0FF3F7FFFFFFFFFFFF),
.INIT_2F(256'hFFFFFFFFFFFFFFF3FFFFFFFFFFF97030FFFFFFFFFFFFFFEFFFFFB130001C1E0E),
.INIT_30(256'h0000000000000000FFFFFFFFFFFFFFF7FFFFFFFFFF9F0E0CFFFFFFFFFFFFFFCF),
.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB({dib[6+0],dib[4+0],dib[2+0],dib[0+0]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+0],dob[4+0],dob[2+0],dob[0+0]}),
      .SSRB(ssrb)
      );

    RAMB16_S1_S4 #(
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h006363F763F763630000000000C6C6C600810081818181810000000000000000),
.INIT_09(256'h00000000000381C000B366D683C6C6830060660381C066060081E7B0E386F3C0),
.INIT_0A(256'h00008181E7818100000081E7C3E78100000381C0C0C0810300C08103030381C0),
.INIT_0B(256'h0000060381C06000008181000000000000000000E70000000381810000000000),
.INIT_0C(256'h00C36660C16066C300E70381C06066C300E781818181838100C36667E7E666C3),
.INIT_0D(256'h0003030381C060E700C36666C70603C100C3666060C706E700C0C0E7C6C3C1C0),
.INIT_0E(256'h038181008181000000818100818100000083C060E36666C300C36666C36666C3),
.INIT_0F(256'h0081008181C066C3000381C060C08103000000E700E7000000C08103060381C0),
.INIT_10(256'h00C36606060666C300C76666C76666C700666666E76666C300C306E6A6E666C3),
.INIT_11(256'h00C36666E60666C300060606C70606E700E70606C70606E70087C6666666C687),
.INIT_12(256'h0066C6870787C6660083C6C0C0C0C0E300E78181818181E700666666E7666666),
.INIT_13(256'h00C36666666666C3006666E6E7676666003636B6B6F7773600E7060606060606),
.INIT_14(256'h00C36660C30666C3006666C6C76666C70063C6A6666666C300060606C76666C7),
.INIT_15(256'h003677F7B6B636360081C3666666666600C366666666666600818181818181E7),
.INIT_16(256'h00C70606060606C700E7060381C060E700818181C3666666006666C381C36666),
.INIT_17(256'hFF00000000000000000000002466C38100E36060606060E3000060C081030600),
.INIT_18(256'h00C3660666C3000000C7666666C7060600E366E360C3000000E70303C70363C1),
.INIT_19(256'hC360E36666E3000000030303C70303C100C306E766C3000000E3666666E36060),
.INIT_1A(256'h0066C687C6660606078181818183008100C38181818300810066666666C70606),
.INIT_1B(256'h00C3666666C300000066666666C700000036B6B6F763000000C3818181818183),
.INIT_1C(256'h00C760C306E300000006060667C600007060E36666E300000606C76666C70000),
.INIT_1D(256'h0063F7B6B63600000081C3666666000000E366666666000000C1030303C70303),
.INIT_1E(256'h00C08181078181C000E70381C0E70000C360E366666600000066C381C3660000),
.INIT_1F(256'hFFFFFFFFFFFFFFFF000000000064B61300038181E08181030081818100818181),
.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_25(256'h7030303030000000000000000000000000000000000000000000000000000000),
.INIT_26(256'hF3F3F7FFFF8F0F06000000001010000000000000000000000E0C0C0C0C000000),
.INIT_27(256'h0000000008080000CFCFEFFFFFF1F060FFFFFFFFFFEF0F0EFFFFFFFFFFF7F070),
.INIT_28(256'h1010103070F0F7FF0808080C0E0FEFFFFFFFFFFFF7F7F3F3F310000000000000),
.INIT_29(256'h0000000000000000C7E1F07030000000CF08000000000000FFFFFFFFEFEFCFCF),
.INIT_2A(256'h000000000000000000000010F0F3F3F3F0F1EFEF8F0000000F8FF7F7F1000000),
.INIT_2B(256'h000000080FCFCFCF000000000000000070303010100000000E0C0C0808000000),
.INIT_2C(256'h1000000000000000F0F0F0F0F0F0F0F000000000000000000000000000000387),
.INIT_2D(256'hF3FFEFCFCFCFCFEF303030707070F0F00C0C0C0E0E0E0F0FCFFFF7F3F3F3F3F7),
.INIT_2E(256'h0000F1F7F78F0F0F000000000000000000000000000000000800000000000000),
.INIT_2F(256'h0000000000000000000000000000068F000000000000000000008FEFEFF1F0F0),
.INIT_30(256'h0000000000000000000000000000000000000000000060F10000000000000000),
.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB({dib[6+1],dib[4+1],dib[2+1],dib[0+1]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+1],dob[4+1],dob[2+1],dob[0+1]}),
      .SSRB(ssrb)
      );
`endif

endmodule


module RAM_PAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );

	 
`ifdef GENERIC_RAM
	wire [15:0] tWire;
	
	sramb16DErsws #(
	.ADDR_WIDTH(10),
	.DATA_WIDTH(16)
	) ram (
		.DIA({DIA,DIA}),
		.WEA(WEA),
		.CLKA(CLKA),
		.ADDRA(ADDRA[10:1]),
		.BEA({ADDRA[0], ~ADDRA[0]}),
		.DOA(tWire),
		
		.DIB(DIB),
		.WEB(WEB),
		.CLKB(CLKB),
		.ADDRB(ADDRB),
		.DOB(DOB)
	);
	
	assign DOA = (ADDRA[0])? tWire[15:8] : tWire[7:0];
	
`else
    RAMB16_S9_S18 #(
      .INIT_00(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_01(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_02(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_03(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_04(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_05(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_06(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_07(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_08(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_09(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_0A(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_0B(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_0C(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_0D(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_0E(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_0F(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_10(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_11(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_12(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_13(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_14(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_15(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_16(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_17(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_18(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_19(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_1A(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_1B(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_1C(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_1D(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_1E(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_1F(256'h7FFF0000000080007FFF0000000080007FFF0000000080007FFF000000008000),.INIT_20(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_21(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_22(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_23(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_24(256'h0000000000008000000000000000800000000000000080000000000000008000),.INIT_25(256'h00002175800010AA00000000800010AA00000000000080000000000000008000),.INIT_26(256'h00002175800010AA00002175800010AA00000000800010AA00002175800010AA),.INIT_27(256'h00002175800010AA00002175800010AA00002175800010AA00002175800010AA),.INIT_28(256'h00002175800010AA00002175800010AA00002175800010AA00002175800010AA),.INIT_29(256'h000000002CA5800020842CA58000184200002175800010AA00002175800010AA),.INIT_2A(256'h00000000217510AA00002175800010AA20842CA58000184220842CA580001842),.INIT_2B(256'h00002175800010AA00000000217510AA00002175800010AA00002175800010AA),.INIT_2C(256'h00002175800010AA00002CA580001842000000002CA5800020842CA580001842),.INIT_2D(256'h00002175800010AA00002175800010AA00002175800010AA00002175800010AA),.INIT_2E(256'h20842CA580001842000000002CA58000000000002CA5800000002175800010AA),.INIT_2F(256'h00000000800010AA00002175800010AA00000000800010AA20842CA580001842),.INIT_30(256'h000000000000000000000000800010AA00002175800010AA00000000800010AA),.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );
`endif

endmodule


module RAM_SPRVAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [31:0] DIB,
    output [31:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [8:0] ADDRB
    );

    RAMB16_S9_S36 #(
      .INIT_00(256'h068C6018067C4018046C601804B7400802A76008029740080087600800774008),.INIT_01(256'h0EA760280E9740280C8760280C7740280A6760280ABC401808AC6018089C4018),.INIT_02(256'h16B7603816A740381497603814874038127760381267403810C7602810B74028),.INIT_03(256'h1E7060581EB940481CA960481C9940481A8960481A7940481869604818C74038),.INIT_04(256'h26A1606826914068248160682471406822B0605822A040582090605820804058),.INIT_05(256'h2E9260882E8240882C7260882CA340782A9360782A8340782873607828B14068),.INIT_06(256'h368E60A8367E40A8346E60A8349E4098328E6098327E4098306E609830A24088),.INIT_07(256'h3E7760C83E6740C83CAD60B83C9D40B83A8D60B83A7D40B8386D60B8389E40A8),.INIT_08(256'h46AB60D8469B40D8448B60D8447B40D8426B60D842A740C8409760C8408740C8),.INIT_09(256'h4E9B60F84E8B40F84C7B60F84C6B40F84A9F60E84A8F40E8487F60E8486F40E8),.INIT_0A(256'h567F6118566F411854AB6108549B4108528B6108527B4108506B610850AB40F8),.INIT_0B(256'h5EAC61285E9C41285C8C61285C7C41285A6C61285AAF4118589F6118588F4118),.INIT_0C(256'h666A614866BC413864AC6138649C4138628C6138627C4138606C613860BC4128),.INIT_0D(256'h6E7A61586E6A41586CCA61486CBA41486AAA61486A9A4148688A6148687A4148),.INIT_0E(256'h76906168768041687470616874CA415872BA615872AA4158709A6158708A4158),.INIT_0F(256'h019001907EAC41787C9C61787C8C41787A7C61787AC0416878B0616878A04168),.INIT_10(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_11(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_12(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_13(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_14(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_15(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_16(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_17(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_18(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_19(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_1A(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_1B(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_1C(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_1D(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_1E(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_1F(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_20(256'h060602500606071007070388070701C40808025A08080138090901220D0D012D),.INIT_21(256'h0404096B050501CE050501B9050507060505071B05050265050504B50606037D),.INIT_22(256'h030303930303096003030976040404C004040E0C040405E3040404AB040400A1),.INIT_23(256'h030312D70303095603030E01030302F1030305D8030312C10303041F03030E16),.INIT_24(256'h02020414020212E202020BC6020212B703031C4D030312CC03031C43030306FB),.INIT_25(256'h020212AC02020E2102020BBB020205EE02022A4402021C380202083302021C22),.INIT_26(256'h02022A6F020202E6020212EC02022583020204290202054C02022A3902020726),.INIT_27(256'h020238860202054102020BB10202037202021C180202083E02021C58020202FC),.INIT_28(256'h0505098C050513380505134D060613430808101008080FF00D0D0FFB0E0E1006),.INIT_29(256'h040409760404135804040664040409810404132D0404101B0404065905050996),.INIT_2A(256'h03030FDB03030CDE04040FD004040CB304040A1704040A22040412EC0404130D),.INIT_2B(256'h0303064E0303122B0303130203030A0D0303132203030CA8030309A1030312F7),.INIT_2C(256'h0303050B0303067A03030CBE0303123503030FE5030312E203030CD303031026),.INIT_2D(256'h02021318020209600202124002020CC902020FC50202066F020209AC02020A2D),.INIT_2E(256'h020213630202033202020CE9020211DF020211D5020212000202108702020516),.INIT_2F(256'h02020644020211CA020210310202095602020F7A02020FA502020A0202020F44),.INIT_30(256'h0606027006060BF106060900070701C40707025A07070BFC080801CE0A0A0265),.INIT_31(256'h040413220404132D05051757050513CF050508F505050C93050513C406061762),.INIT_32(256'h0303090A03030F9A0303018E03030C070404176C04040199040401D904040C9D),.INIT_33(256'h03030FA503030F8F030304CB03030D29030313B90303119403031E9303031189),.INIT_34(256'h030305F803030D3403030869030315880303159303031E8803030ACF03031031),.INIT_35(256'h0202119F0202013802020C88020228B60202117E020205620202174C02020AC4),.INIT_36(256'h020210260202039302021A5E0202012D02021A5302020B2F02021798020204D6),.INIT_37(256'h02021F1F0202033D020228AB0202178D0202039D0202120002021AF502020F84),.INIT_38(256'h6620313130322031323A37323A36302035322079614D2064655720746C697542),.INIT_39(256'h202020202020202020202020202020204D3239393A393839206E7673206D6F72),.INIT_3A(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_3B(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_3C(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_3D(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_3E(256'h0190019001900190019001900190019001900190019001900190019001900190),.INIT_3F(256'h0190019001900190019001900190019001900190019001900190019001900190)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_SPRPAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );
`ifdef GENERIC_RAM
	wire [15:0] tWire;
	
	sramb16DErsws #(
	.ADDR_WIDTH(10),
	.DATA_WIDTH(16)
	) ram (
		.DIA({DIA,DIA}),
		.WEA(WEA),
		.CLKA(CLKA),
		.ADDRA(ADDRA[10:1]),
		.BEA({ADDRA[0], ~ADDRA[0]}),
		.DOA(tWire),
		
		.DIB(DIB),
		.WEB(WEB),
		.CLKB(CLKB),
		.ADDRB(ADDRB),
		.DOB(DOB)
	);
	
	assign DOA = (ADDRA[0])? tWire[15:8] : tWire[7:0];
	
`else
    RAMB16_S9_S18 #(
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_12(256'h0000000000000000000000000000000000000000000000000000000004200421),.INIT_13(256'h0000000000000000000000000000000000000000000000000000002004200421),.INIT_14(256'h0000000000000000000000000000000000000000000000210020042004210421),.INIT_15(256'h0000000000000000000000000000000000000000000000210021042104210421),.INIT_16(256'h0000000000000000000000000000000000000000002100210021042104210421),.INIT_17(256'h0000000000000000000000000000000000000000002100210421042104210842),.INIT_18(256'h0000000000000000000000000000000000000021002100210421044108410842),.INIT_19(256'h0000000000000000000000000000000000000021002104210421044108410842),.INIT_1A(256'h0000000000000000000000000000040104210421042104420441084108420C63),.INIT_1B(256'h0000000000000000000000000000040104210421042104420441084108420C63),.INIT_1C(256'h000000000000000000000000000104210421042104210442044208620C620C63),.INIT_1D(256'h000000000000000000000001040104210421042104420442044208620C620C63),.INIT_1E(256'h000000000000000000000001042104210421042104420442086208620C631084),.INIT_1F(256'h00000000000000000000000104210421042104420442046308620C6210831084),.INIT_20(256'h00000000000000000001040104210421042104420442086308630C83108314A5),.INIT_21(256'h00000000000000000001040104210421084208420842086308830C8314A414A5),.INIT_22(256'h0000000000000000000104210421082208420842086308840C8310A314A418C6),.INIT_23(256'h0000000000000000000104210421082208420842086308840C8310A314A418C6),.INIT_24(256'h0000000000000000000104210422084208420863086308840CA410A418C51CE7),.INIT_25(256'h040000000000000104210422082208420842086308840CA50CA414C418C51CE7),.INIT_26(256'h040000000000000104210422082208420842086308840CA510A414C41CE52108),.INIT_27(256'h040000000000000104210422084208420C630C630C840CA510C514E51CE62108),.INIT_28(256'h04000000000000010421042208420C430C630C630C840CC610C518E521062529),.INIT_29(256'h04000000000000010421042208420C430C630C840CA50CC610E5190521072529),.INIT_2A(256'h04000000000004210422082208430C630C630C840CA510C614E619062527294A),.INIT_2B(256'h04000000000004210422082208430C631084108410A510E715061D2629482D6B),.INIT_2C(256'h0400000000000421042208230C430C63108410A510C610E715071D2729482D6B),.INIT_2D(256'h0400000000000421042208430C431064108410A510C61508192721472D69318C),.INIT_2E(256'h0400000000000421042208430C631064108410A510E71508192721672D6935AD),.INIT_2F(256'h0400000000000421042208430C64108414A514C614E715291D482568318A39CE),.INIT_30(256'h0400000000000421042208430C64108414A514C614E715291D48258835AA39CE),.INIT_31(256'h080000000421042208430C441064148514A514C61508194A1D6929A939CB3DEF),.INIT_32(256'h080000000421042208430C441064148518C618E71908194A218929A939CC4210),.INIT_33(256'h080000000421042208430C44108514A518C618E71929196B218A2DCA3DEC4631),.INIT_34(256'h080000000421042208430C64108518A618C618E719291D8C25AA31EA420D4A52),.INIT_35(256'h080000000421042208430C65148518A61CE71D081D4A1D8C25CB31EB462E4E73),.INIT_36(256'h080000000421084208441065148618C61CE71D081D4A21AD29CC360C4A4E5294),.INIT_37(256'h08000000042108420844106514861CC71CE71D291D6B21CE29EC3A2C4A4F56B5),.INIT_38(256'h08000000042108420844106514A61CC721082129216B21CE2E0D3A4D4E705AD6),.INIT_39(256'h0C000000042108430C64106618A61CC72108214A218C25EF2E0D3E6D52905EF7),.INIT_3A(256'h0C000000042108430C64108618A720E82108214A218C2610322E428E56B16318),.INIT_3B(256'h0C000000042108430C65148618A720E82529254A25AD2A10324F42AF5AD26739),.INIT_3C(256'h0C000000042108430C6514871CC720E82529256B25CE2A31366F46CF5EF36B5A),.INIT_3D(256'h0C000000042108430C6514871CC82509294A296B29CE2E5236904AD063146F7B),.INIT_3E(256'h0C000000042108430C6514871CC82509294A298C29EF2E733AB14EF16735739C),.INIT_3F(256'h1000000008420C64108614A820E9292A2D6B2DAD2E1032943ED253326F767BDE)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );
`endif

endmodule


module RAM_CODEL (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
`ifdef ALTERA
  output [7:0] ao,
  output [7:0] bo
`else
   output reg [7:0] ao,
  output reg [7:0] bo
`endif
  );

  
`ifdef GENERIC_RAM
	srambDrsws #(
		.DATA_WIDTH(8),
		.ADDR_WIDTH(7)
	) ram (
		.DIA(ad),
      .WEA(wea),
      .CLKA(wclk),
      .ADDRA(a),
      .DOA(ao),

      .DIB(8'b00000000),
      .WEB(0),
      .CLKB(wclk),
      .ADDRB(b),
      .DOB(bo),
	);
	
`elsif ALTERA
	// NOTE: This does not have a clocked output register
	RAM128X8D ram(
        .D(ad),
        .WE(wea),
        .WCLK(wclk),
        .A(a),
        .DPRA(b),
        .SPO(ao),
        .DPO(bo)
		  );

`else

  wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end
      mRAM128X1D
      #( .INIT(128'b00101101010101011110101000110001000101010111110101010010010111110100000101111001001011010001101000101111100101100100000111110010) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
      #( .INIT(128'b11100001010110100111100000010010000100110011101101000010001011110001010010100001101101010000000001000011100101000101101010110011) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
      #( .INIT(128'b01010001011010001100010000010000111000000010101000000000011010000101011000100000100100000110000111000100100001001100100010101000) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
      #( .INIT(128'b10100000000100010100000000100001100000000000100000000000010010000100000000000001110100000100000000000100100001010100000010101001) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
      #( .INIT(128'b10100000000100000000000000000001000000000000101000000010000000010000000000000001000100000000000000000000100001000000000000000000) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
      #( .INIT(128'b10000100010000010000000000000100000000000010100000000010000100010000000000000100000000001010100000000000100001000000000000010000) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
      #( .INIT(128'b10000001011000111000000000010100110000000000001000100000000000000000000000110010000000000000000000000000100001001000000000000001) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
      #( .INIT(128'b11101101011101111100001000010111111001100110011010110010011100010111111111011001010010000011101111101100101001110001111100000001) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));
`endif

endmodule


module RAM_CODEH (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
`ifdef ALTERA
  output [7:0] ao,
  output [7:0] bo
`else
   output reg [7:0] ao,
  output reg [7:0] bo
`endif
  );


`ifdef GENERIC_RAM
	srambDrsws #(
		.DATA_WIDTH(8),
		.ADDR_WIDTH(7)
	) ram (
		.DIA(ad),
      .WEA(wea),
      .CLKA(wclk),
      .ADDRA(a),
      .DOA(ao),

      .DIB(8'b00000000),
      .WEB(0),
      .CLKB(wclk),
      .ADDRB(b),
      .DOB(bo),
	);
	
`elsif ALTERA
	// NOTE: This does not have a clocked output register
	RAM128X8D ram(
        .D(ad),
        .WE(wea),
        .WCLK(wclk),
        .A(a),
        .DPRA(b),
        .SPO(ao),
        .DPO(bo)
		  );

`else
    wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end
      mRAM128X1D
      #( .INIT(128'b11100101011100111100100010111110111001100011001101000111011111110111111111110001010000010011101111101101101101010001111000100001) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
      #( .INIT(128'b00000000100000000010000000000000000110010001000101000000110000001100000000000000001001000000010000010101010110000010000010000000) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
      #( .INIT(128'b11100101111100111100100000011110111000101010001100000010011100010001011010010001010000010011101111010010000010010111101000001001) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
      #( .INIT(128'b00010000000010000000100000000001000010000000000000000000100000001100000000000010100000110000010000010100010000000010000000001010) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
      #( .INIT(128'b11100101111100111101000000011110111000101010001000000010011110010001011010010001010000100111101111000000000000010101101010101001) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
      #( .INIT(128'b00011000110011010011101000001101100111011101011101010000110011101110100101111010101011110110110000111111011110101110010110111110) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
      #( .INIT(128'b01101101001101101110101000010010011101110111010101010000011111101111111111101001011011010101011011111111011110111111111110111100) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
      #( .INIT(128'b00010010100010000001010111101001000010001000100010101101100000000000000000000110100100101000000000000000100001000000000001000010) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));
`endif
endmodule

