
module RAM_SPRIMG (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [14:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [14:0] addrb
    );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB(dib[0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[0]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB(dib[1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[1]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram2 (
      .DIA(dia[2]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[2]),
      .SSRA(ssra),

      .DIB(dib[2]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[2]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram3 (
      .DIA(dia[3]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[3]),
      .SSRA(ssra),

      .DIB(dib[3]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[3]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
      .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram4 (
      .DIA(dia[4]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4]),
      .SSRA(ssra),

      .DIB(dib[4]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram5 (
      .DIA(dia[5]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[5]),
      .SSRA(ssra),

      .DIB(dib[5]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[5]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
         .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram6 (
      .DIA(dia[6]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[6]),
      .SSRA(ssra),

      .DIB(dib[6]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[6]),
      .SSRB(ssrb)
      );

    RAMB16_S1_S1 #(
            .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram7 (
      .DIA(dia[7]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[7]),
      .SSRA(ssra),

      .DIB(dib[7]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[7]),
      .SSRB(ssrb)
      );

endmodule


module RAM_PICTURE (
    input [7:0] dia,
    output [7:0] doa,
    input wea,
    input ena,
    input clka,
    input ssra,
    input [12:0] addra,
    input [7:0] dib,
    output [7:0] dob,
    input web,
    input enb,
    input clkb,
    input ssrb,
    input [12:0] addrb
    );

    RAMB16_S4_S4 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram0 (
      .DIA(dia[4*0+3:4*0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*0+3:4*0]),
      .SSRA(ssra),

      .DIB(dib[4*0+3:4*0]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*0+3:4*0]),
      .SSRB(ssrb)
      );

    RAMB16_S4_S4 #(
          .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram1 (
      .DIA(dia[4*1+3:4*1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[4*1+3:4*1]),
      .SSRA(ssra),

      .DIB(dib[4*1+3:4*1]),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB(dob[4*1+3:4*1]),
      .SSRB(ssrb)
      );

endmodule


module RAM_CHR (
    input [1:0] dia, 	// NC
    output [1:0] doa, 	// CHAROUT
    input wea, 		// 0
    input ena,   	// 1
    input clka,		// vga_clk
    input ssra,		// 0
    input [14:0] addra,	// {glyph, row[2:0], _column[2], ~_column[1:0]}
    input [7:0] dib,	// mem_data_wr
    output [7:0] dob,	// mem_data_rd1
    input web,		// mem_wr
    input enb,		// en_chr
    input clkb,		// mem_clk
    input ssrb,		// 0
    input [12:0] addrb	// mem_addr
    );

// 32 across
// Address mode:  AAAAAA / B BBBB, where A is the INIT_A, and B is the bit across the line
//      Note bit 255 .... bit 0
// Note that ASCII 64, hex 0x40 starts at address 0x0400 
    RAMB16_S1_S4 #(
.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
// Hex 0x20 below
.INIT_08(256'h006666FF66FF6666_0000000000666666_0081000081818181_0000000000000000),
.INIT_09(256'h000000000081C060_00F3667683C366C3_0064660381C06626_0081C760C306E381),
.INIT_0A(256'h00008181E7818100_000066C3FFC36600_000381C0C0C08103_00C08103030381C0),
.INIT_0B(256'h00060381C0603000_0081810000000000_00000000E7000000_0381810000000000),
.INIT_0C(256'h00C36660C16066C3_00E70603C06066C3_00E7818181838181_00C3666667E666C3),
.INIT_0D(256'h0081818181C066E7_00C36666C70666C3_00C3666060C706E7_006060F766E1E060),
.INIT_0E(256'h0381810000810000_0000810000810000_00C36660E36666C3_00C36666C36666C3),
.INIT_0F(256'h00810081C06066C3_000781C060C08107_000000E700E70000_00E08103060381E0),
//       Character 0x40 starts on the line below
.INIT_10(256'h00C36606060666C3_00C76666C76666C7_00666666E766C381_00C32606E6E666C3),
.INIT_11(256'h00C36666E60666C3_00060606870606E7_00E70606870606E7_0087C6666666C687),
.INIT_12(256'h0066C6870787C666_0083C6C0C0C0C0E1_00C38181818181C3_00666666E7666666),
.INIT_13(256'h00C36666666666C3_006666E6E7E76766_00363636B6F77736_00E7060606060606),
.INIT_14(256'h00C36660C30666C3_0066C687C76666C7_00E0C366666666C3_00060606C76666C7),
.INIT_15(256'h003677F7B6363636_0081C36666666666_00C3666666666666_00818181818181E7),
.INIT_16(256'h00C30303030303C3_00E7060381C060E7_00818181C3666666_006666C381C36666),
.INIT_17(256'h00E7000000000000_0000000066C38100_00C3C0C0C0C0C0C3_003060C081030600),
.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram0 (
      .DIA(dia[0]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[0]),
      .SSRA(ssra),

      .DIB({dib[6+0],dib[4+0],dib[2+0],dib[0+0]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+0],dob[4+0],dob[2+0],dob[0+0]}),
      .SSRB(ssrb)
      );

    // note: for [A | B] 6C produces [B | A]

    RAMB16_S1_S4 #(
.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
// hex 0x20 below
.INIT_08(256'h006666FF66FF6666_0000000000666666_0081000081818181_0000000000000000),
.INIT_09(256'h000000000081C060_00F3667683C366C3_0064660381C06626_0081C760C306E381),
.INIT_0A(256'h00008181E7818100_000066C3FFC36600_000381C0C0C08103_00C08103030381C0),
.INIT_0B(256'h00060381C0603000_0081810000000000_00000000E7000000_0381810000000000),
.INIT_0C(256'h00C36660C16066C3_00E70603C06066C3_00E7818181838181_00C3666667E666C3),
.INIT_0D(256'h0081818181C066E7_00C36666C70666C3_00C3666060C706E7_006060F766E1E060),
.INIT_0E(256'h0381810000810000_0000810000810000_00C36660E36666C3_00C36666C36666C3),
.INIT_0F(256'h00810081C06066C3_000781C060C08107_000000E700E70000_00E08103060381E0),
//       Character 0x40 starts on the line below
.INIT_10(256'h00C36606060666C3_00C76666C76666C7_00666666E766C381_00C32606E6E666C3),
.INIT_11(256'h00C36666E60666C3_00060606870606E7_00E70606870606E7_0087C6666666C687),
.INIT_12(256'h0066C6870787C666_0083C6C0C0C0C0E1_00C38181818181C3_00666666E7666666),
.INIT_13(256'h00C36666666666C3_006666E6E7E76766_00363636B6F77736_00E7060606060606),
.INIT_14(256'h00C36660C30666C3_0066C687C76666C7_00E0C366666666C3_00060606C76666C7),
.INIT_15(256'h003677F7B6363636_0081C36666666666_00C3666666666666_00818181818181E7),
.INIT_16(256'h00C30303030303C3_00E7060381C060E7_00818181C3666666_006666C381C36666),
.INIT_17(256'h00E7000000000000_0000000066C38100_00C3C0C0C0C0C0C3_003060C081030600),
.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram1 (
      .DIA(dia[1]),
      .WEA(wea),
      .ENA(ena),
      .CLKA(clka),
      .ADDRA(addra),
      .DOA(doa[1]),
      .SSRA(ssra),

      .DIB({dib[6+1],dib[4+1],dib[2+1],dib[0+1]}),
      .WEB(web),
      .ENB(enb),
      .CLKB(clkb),
      .ADDRB(addrb),
      .DOB({dob[6+1],dob[4+1],dob[2+1],dob[0+1]}),
      .SSRB(ssrb)
      );

endmodule


module RAM_PAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );

    RAMB16_S9_S18 #(
      	.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_SPRVAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [31:0] DIB,
    output [31:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [8:0] ADDRB
    );

    RAMB16_S9_S36 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_SPRPAL (
    input [7:0] DIA,
    output [7:0] DOA,
    input WEA,
    input ENA,
    input CLKA,
    input SSRA,
    input [10:0] ADDRA,
    input [15:0] DIB,
    output [15:0] DOB,
    input WEB,
    input ENB,
    input CLKB,
    input SSRB,
    input [9:0] ADDRB
    );

    RAMB16_S9_S18 #(
           .INIT_00(0),
.INIT_01(0),
.INIT_02(0),
.INIT_03(0),
.INIT_04(0),
.INIT_05(0),
.INIT_06(0),
.INIT_07(0),
.INIT_08(0),
.INIT_09(0),
.INIT_0A(0),
.INIT_0B(0),
.INIT_0C(0),
.INIT_0D(0),
.INIT_0E(0),
.INIT_0F(0),
.INIT_10(0),
.INIT_11(0),
.INIT_12(0),
.INIT_13(0),
.INIT_14(0),
.INIT_15(0),
.INIT_16(0),
.INIT_17(0),
.INIT_18(0),
.INIT_19(0),
.INIT_1A(0),
.INIT_1B(0),
.INIT_1C(0),
.INIT_1D(0),
.INIT_1E(0),
.INIT_1F(0),
.INIT_20(0),
.INIT_21(0),
.INIT_22(0),
.INIT_23(0),
.INIT_24(0),
.INIT_25(0),
.INIT_26(0),
.INIT_27(0),
.INIT_28(0),
.INIT_29(0),
.INIT_2A(0),
.INIT_2B(0),
.INIT_2C(0),
.INIT_2D(0),
.INIT_2E(0),
.INIT_2F(0),
.INIT_30(0),
.INIT_31(0),
.INIT_32(0),
.INIT_33(0),
.INIT_34(0),
.INIT_35(0),
.INIT_36(0),
.INIT_37(0),
.INIT_38(0),
.INIT_39(0),
.INIT_3A(0),
.INIT_3B(0),
.INIT_3C(0),
.INIT_3D(0),
.INIT_3E(0),
.INIT_3F(0)
    ) ram (
      .DIPA(0),
      .DIA(DIA),
      .WEA(WEA),
      .ENA(ENA),
      .CLKA(CLKA),
      .ADDRA(ADDRA),
      .DOA(DOA),
      .SSRA(SSRA),

      .DIPB(0),
      .DIB(DIB),
      .WEB(WEB),
      .ENB(ENB),
      .CLKB(CLKB),
      .ADDRB(ADDRB),
      .DOB(DOB),
      .SSRB(SSRB)
      );

endmodule


module RAM_CODEL (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
  output reg [7:0] ao,
  output reg [7:0] bo
  );
  wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end

      mRAM128X1D
      #( .INIT(0) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
      #( .INIT(0) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
      #( .INIT(0) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
      #( .INIT(0) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
      #( .INIT(0) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
      #( .INIT(0) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
      #( .INIT(0) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
      #( .INIT(0) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));

endmodule


module RAM_CODEH (
  input wclk,
  input [7:0] ad,
  input wea,
  input [6:0] a,
  input [6:0] b,
  output reg [7:0] ao,
  output reg [7:0] bo
  );
  wire [7:0] _ao;
  wire [7:0] _bo;
  always @(posedge wclk)
  begin
    ao <= _ao;
    bo <= _bo;
  end

      mRAM128X1D
           #( .INIT(0) )
      ram0(
        .D(ad[0]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[0]),
        .DPO(_bo[0]));

      mRAM128X1D
           #( .INIT(0) )
      ram1(
        .D(ad[1]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[1]),
        .DPO(_bo[1]));

      mRAM128X1D
           #( .INIT(0) )
      ram2(
        .D(ad[2]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[2]),
        .DPO(_bo[2]));

      mRAM128X1D
           #( .INIT(0) )
      ram3(
        .D(ad[3]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[3]),
        .DPO(_bo[3]));

      mRAM128X1D
           #( .INIT(0) )
      ram4(
        .D(ad[4]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[4]),
        .DPO(_bo[4]));

      mRAM128X1D
            #( .INIT(0) )
      ram5(
        .D(ad[5]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[5]),
        .DPO(_bo[5]));

      mRAM128X1D
          #( .INIT(0) )
      ram6(
        .D(ad[6]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[6]),
        .DPO(_bo[6]));

      mRAM128X1D
            #( .INIT(0) )
      ram7(
        .D(ad[7]),
        .WE(wea),
        .WCLK(wclk),
        .A0(a[0]),
        .A1(a[1]),
        .A2(a[2]),
        .A3(a[3]),
        .A4(a[4]),
        .A5(a[5]),
        .A6(a[6]),
        .DPRA0(b[0]),
        .DPRA1(b[1]),
        .DPRA2(b[2]),
        .DPRA3(b[3]),
        .DPRA4(b[4]),
        .DPRA5(b[5]),
        .DPRA6(b[6]),
        .SPO(_ao[7]),
        .DPO(_bo[7]));

endmodule

